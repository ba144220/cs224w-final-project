module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;

    assign temp_0 = $signed(($unsigned(($signed(($unsigned(($unsigned(input_data) * input_data)) * input_data)) & input_data)) * input_data));
    assign temp_1 = temp_0 ? ($signed(($signed(($signed(($signed(($signed(($unsigned(($unsigned(($unsigned((($signed(($signed(temp_0) & temp_0)) + temp_0) & temp_0)) * temp_0[6:6])) + temp_0)) | temp_0)) & input_data)) | (~temp_0))) | temp_0)) - (~temp_0))) * temp_0) : ($signed(($signed(($unsigned(($unsigned(($signed(($signed(($unsigned(($unsigned(($signed(temp_0[6:2]) | input_data)) * temp_0)) + input_data)) * temp_0)) & temp_0[6:5])) & input_data)) | temp_0)) | input_data)) + temp_0[6:5]);
    logic [31:0] expr_86570;
    assign expr_86570 = ($unsigned((($signed(($signed(($signed(($unsigned(temp_1) ^ temp_0)) + temp_0)) * temp_0[6:3])) | temp_0) ^ temp_0)) | temp_1);
    assign temp_2 = expr_86570[30:0];
    assign temp_3 = (($unsigned((($unsigned(($unsigned(($signed(($unsigned(($unsigned(($unsigned((input_data ^ temp_0)) * temp_1)) * temp_0)) + temp_1)) ^ temp_2)) | temp_1)) & temp_1) & temp_0)) * temp_1) | temp_0[6:2]);
    assign temp_4 = ($signed(($unsigned((($signed(($signed(($signed(($unsigned(($unsigned(temp_0) + temp_0)) - temp_1)) | temp_3)) * (~temp_2))) ^ temp_1[25:20]) & input_data)) ^ input_data)) | input_data);
    logic [10:0] expr_377313;
    assign expr_377313 = $signed(($signed(($unsigned(($signed((temp_0 + temp_0)) + temp_0)) + temp_4)) | temp_0));
    assign temp_5 = expr_377313[4:0];
    assign temp_6 = ($unsigned(($unsigned(($unsigned(($unsigned(($unsigned(($unsigned(((($unsigned(($unsigned(($unsigned(temp_3) - temp_0)) ^ temp_2[30:29])) & input_data[4:3]) | temp_3) * temp_1)) - temp_3)) + temp_0)) ^ temp_1)) * temp_2)) - (~temp_1[25:6]))) * temp_5);
    assign temp_7 = ($signed(($signed(($signed(($unsigned(($unsigned(($signed(temp_0) * temp_4)) + (~input_data))) + temp_6)) ^ temp_1)) - temp_5)) | temp_0);
    assign temp_8 = temp_0;
    assign temp_9 = $signed(($signed(($signed(((($unsigned(temp_8) * temp_5[4:2]) & temp_1) ^ temp_0)) + temp_2)) - temp_4));
    assign temp_10 = ($signed(($unsigned(($signed(($signed(($unsigned(temp_6[1:1]) ^ input_data)) + temp_0)) * temp_3)) - temp_8)) ^ temp_9[3:2]);
    assign temp_11 = $signed(($signed(($unsigned(($unsigned(($unsigned(($unsigned(($signed((($unsigned(temp_7) + temp_9) ^ temp_5)) ^ temp_7)) - temp_5)) | temp_0)) ^ temp_3)) + (~temp_0))) - input_data));
    assign temp_12 = ($unsigned((($unsigned(($signed(($unsigned(($signed(($unsigned((($unsigned(temp_1) + temp_1) * temp_4)) * temp_8)) | temp_2)) ^ temp_10)) & temp_8[18:1])) ^ temp_3) ^ temp_7)) ^ temp_9);
    assign temp_13 = ($unsigned(($unsigned(temp_7) * temp_0)) | temp_12[17:15]);

    logic [20:0] expr_817517;
    assign expr_817517 = ($signed(($unsigned(temp_3) + temp_8)) ^ temp_10[14:5]);
    assign output_data = expr_817517[19:0];

endmodule