module top (
    input [7:0] input_data,
    output [9:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;
    logic [26:0] temp_10;
    logic [4:0] temp_11;
    logic [15:0] temp_12;
    logic [5:0] temp_13;
    logic [27:0] temp_14;
    logic [3:0] temp_15;
    logic [7:0] temp_16;
    logic [14:0] temp_17;

    assign temp_0 = ((((input_data + input_data) + input_data) - input_data) & input_data);
    assign temp_1 = (temp_0 * temp_0[14:0]);
    assign temp_2 = input_data[6:2];
    assign temp_3 = (((temp_2[4:3] == temp_2) + input_data[6:0]) | temp_0);
    assign temp_4 = (((temp_2 - temp_1[3:0]) | temp_2[4:0]) * input_data);
    assign temp_5 = (((temp_0 & temp_2) * temp_0) * temp_3[4:0]);
    assign temp_6 = ((temp_4[17:0] * temp_4) + temp_2);
    assign temp_7 = $signed(((((temp_6 - temp_3[6:1]) - temp_2) * temp_0) | temp_3));
    assign temp_8 = (temp_6 + temp_2[4:4]);
    assign temp_9 = (($signed(temp_1) < input_data) >= temp_8);
    assign temp_10 = (((temp_2[4:4] - temp_2[4:0]) + temp_8) + temp_4[4:0]);
    assign temp_11 = ((((temp_4 & temp_3) | temp_3) + temp_6[11:0]) - input_data[6:2]);
    assign temp_12 = (((temp_3[4:0] | temp_6) | temp_11[3:0]) + temp_3);
    assign temp_13 = $unsigned((($unsigned((input_data[7:2] | temp_11)) + temp_0) + temp_5));
    assign temp_14 = ((temp_4 > temp_2) + temp_8);
    assign temp_15 = ((((temp_11 - temp_11) - temp_10) & temp_10) - temp_7[2:0]);
    assign temp_16 = ((temp_2 - temp_0[3:0]) & temp_9[27:17]);
    assign temp_17 = $unsigned(((temp_4[23:0] | temp_16[5:0]) + temp_7[1:0]));

    assign output_data = ((((temp_0[25:17] | temp_2[4:4]) * temp_7) & temp_12[15:0]) | temp_6[3:0]);

endmodule