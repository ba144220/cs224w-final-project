module top (
    input [5:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;

    assign temp_0 = $unsigned((25'd27357858 & input_data));
    assign temp_1 = input_data;
    assign temp_2 = input_data[1:1] ? input_data : ($unsigned(temp_1) & temp_0);
    assign temp_3 = ($signed(temp_1[5:0]) << temp_2);
    assign temp_4 = ($unsigned(temp_1) - (~temp_3));
    assign temp_5 = $unsigned(input_data);
    assign temp_6 = $unsigned(16'd27535);
    assign temp_7 = $signed(($unsigned(($unsigned(temp_0[20:0]) - temp_3)) ^ temp_5[8:0]));
    assign temp_8 = temp_5;
    assign temp_9 = ($unsigned((temp_6 + temp_4)) - temp_1);
    assign temp_10 = (temp_6 | temp_6);
    assign temp_11 = (temp_8 + temp_4);
    assign temp_12 = {20'b0, $signed(($signed(temp_5) | temp_3))};
    assign temp_13 = ($signed((temp_2[4:0] ^ temp_1)) + temp_5);
    assign temp_14 = {23'b0, temp_5};

    assign output_data = ($unsigned(($signed(temp_2) & temp_11)) ^ temp_3);

endmodule