module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;
    logic [17:0] temp_12;
    logic [2:0] temp_13;
    logic [1:0] temp_14;
    logic [23:0] temp_15;
    logic [29:0] temp_16;
    logic [20:0] temp_17;

    assign temp_0 = ($signed(($signed(($signed(($unsigned(($unsigned(($signed(input_data) - 6'd17)) | input_data)) * input_data)) & input_data)) & input_data)) * input_data);
    assign temp_1 = {14'b0, $unsigned(($signed(((($unsigned(temp_0) | temp_0) + temp_0) | temp_0)) ^ temp_0))};
    assign temp_2 = ($signed(($unsigned(temp_0) + temp_0)) + input_data);
    assign temp_3 = $signed(($unsigned((temp_1 * temp_1)) * temp_0));
    assign temp_4 = temp_1 ? ($signed(((($unsigned(($signed(temp_0) - temp_0[5:2])) ^ temp_2) & temp_0[5:4]) + temp_3)) * temp_2) : (($signed((($signed(($signed(($unsigned(($signed(temp_0[1:0]) * temp_0)) - temp_3)) & input_data)) ^ temp_2) ^ input_data)) - temp_2) | temp_2);
    assign temp_5 = ($unsigned(($signed(($unsigned(($unsigned(($unsigned(($signed((($signed(($unsigned(($signed(temp_2) + temp_3)) & input_data)) & temp_4) * temp_3)) ^ input_data)) & input_data)) & temp_0[2:0])) + temp_4)) | temp_4)) + temp_3);
    assign temp_6 = ($signed(($signed((($unsigned(($signed(($signed(($signed(temp_1) & temp_5)) & temp_1[18:0])) & temp_1)) * temp_2) + temp_1)) ^ temp_0)) + temp_3);
    assign temp_7 = ($unsigned(($signed(temp_2[10:4]) & temp_5)) | temp_3);
    assign temp_8 = $signed((($signed(($unsigned(($unsigned((($unsigned(input_data) | temp_1) & temp_2)) - temp_6[2:0])) * temp_2)) * temp_6[2:1]) * input_data));
    assign temp_9 = ($unsigned(($unsigned(($signed((($signed(($signed(($signed(($signed(($unsigned(temp_6[2:2]) & temp_5)) & input_data)) + temp_2)) & temp_0)) + temp_7) - temp_8)) | temp_8)) + temp_0)) ^ temp_2);
    assign temp_10 = ($unsigned(($unsigned(temp_8) | temp_4)) | temp_3);
    assign temp_11 = temp_3 ? $unsigned(temp_8) : ($unsigned(($signed(($signed(($unsigned((($unsigned(($signed(($signed(($signed(($signed(temp_4) + temp_6[2:2])) * 29'd280757811)) - temp_2)) & temp_9)) * temp_5) - temp_4)) + temp_5)) + temp_0)) ^ temp_9)) - temp_4);
    assign temp_12 = ($signed(($unsigned(($signed(($signed(($unsigned(($unsigned(temp_10) ^ temp_6)) - temp_8)) & temp_6)) & temp_11)) ^ temp_5[13:3])) | temp_10);
    logic [30:0] expr_244691;
    assign expr_244691 = ($unsigned(($signed(($signed(((temp_9 ^ temp_7) * temp_10[22:0])) + temp_1)) - temp_0[3:0])) + input_data);
    assign temp_13 = expr_244691[2:0];
    assign temp_14 = {1'b0, ($signed(temp_4) <= temp_8)};
    assign temp_15 = ($signed(($signed(temp_13) - temp_2)) & temp_4);
    assign temp_16 = temp_0 ? temp_8 : $signed(($signed(($unsigned(($signed(($signed(($signed(((temp_5 * temp_7) | temp_14)) ^ temp_11)) - temp_15)) & temp_8)) + temp_11)) + temp_15));
    assign temp_17 = temp_15 ? temp_7 : ($unsigned(($signed(($unsigned(($unsigned(($unsigned(($unsigned(temp_8) * temp_11)) - temp_14)) & temp_11)) & temp_4)) ^ temp_5)) + temp_15[23:15]);

    logic [32:0] expr_315260;
    assign expr_315260 = (($signed(($unsigned(($signed(($unsigned(((($unsigned(temp_0) + temp_13) ^ temp_10[23:8]) * temp_3)) + temp_8)) ^ temp_4)) + temp_0)) ^ temp_15) ^ temp_4[16:3]);
    logic [36:0] expr_454962;
    assign expr_454962 = $signed(($signed((($signed(($signed(($signed(($signed(($unsigned(($signed((temp_4 | temp_7)) - temp_13[2:2])) - temp_16)) & temp_7)) | temp_5)) - temp_16)) + temp_11[28:4]) * temp_13)) - temp_12[17:10]));
    assign output_data = temp_4 ? expr_315260[5:0] : expr_454962[5:0];

endmodule