module top (
    input [7:0] input_data,
    output [4:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;

    assign temp_0 = input_data[3:3] ? input_data : input_data;
    logic [27:0] expr_585184;
    assign expr_585184 = ((($signed(($signed(input_data[7:4]) >= temp_0[23:0])) == temp_0) & temp_0) - temp_0);
    assign temp_1 = expr_585184[3:0];
    assign temp_2 = (($unsigned(temp_1[1:0]) * temp_0[23:0]) & temp_1);
    assign temp_3 = ($unsigned(($signed(temp_1[2:0]) < temp_0)) < (~input_data[6:0]));
    assign temp_4 = (temp_1 | temp_0);
    assign temp_5 = ($unsigned(((temp_1[3:3] + temp_4[23:12]) & temp_1)) - temp_3);
    assign temp_6 = (temp_4 * input_data);
    assign temp_7 = $unsigned((($signed(((temp_6 & temp_1) * temp_1)) * temp_2[1:0]) | temp_4));

    assign output_data = $signed((temp_5[3:0] & temp_7));

endmodule