module top (
    input [2:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;
    logic [25:0] temp_16;
    logic [5:0] temp_17;

    assign temp_0 = input_data;
    assign temp_1 = $unsigned((temp_0 & (~input_data)));
    assign temp_2 = $signed((($unsigned((((((((temp_1 - input_data) & temp_0) | (~input_data)) * temp_0) - input_data) * temp_1) & (~temp_1))) + input_data) - -13'd576));
    assign temp_3 = $signed((((((((temp_2[6:0] & temp_0) & temp_2) + input_data) + temp_1[4:0]) | input_data) ^ input_data) & input_data));
    assign temp_4 = {5'b0, ((((input_data <= temp_2) ^ temp_2) <= input_data) <= temp_0)};
    assign temp_5 = $unsigned(((((input_data - temp_1) | temp_1) ^ (~temp_4)) | temp_2[8:0]));
    assign temp_6 = {12'b0, (input_data - input_data)};
    assign temp_7 = $signed(((($unsigned(((((((temp_3[1:0] + (~temp_0)) + temp_6) - temp_3[1:0]) - (~temp_1)) & temp_4) ^ input_data)) | temp_2) | temp_4) & temp_0));
    assign temp_8 = temp_2;
    assign temp_9 = $unsigned((((($signed((temp_5 ^ temp_7)) ^ temp_6) ^ (~temp_3)) * temp_0) | temp_7));
    assign temp_10 = $signed((($unsigned((($signed((((($signed((temp_3 - temp_8)) - (~temp_6)) ^ temp_5) | temp_4[2:0]) & temp_0)) ^ temp_6) ^ temp_9)) + temp_7) * temp_9[1:0]));
    assign temp_11 = ((($signed(((($signed((temp_1 | temp_7)) & temp_8) ^ (~temp_3)) * input_data)) + input_data) ^ temp_6) - temp_0);
    assign temp_12 = $signed((($signed((((((((temp_1 - (~temp_5)) >> temp_4) >> temp_3) << input_data) * input_data) * temp_11) << temp_4[2:0])) >> temp_11) - temp_1));
    assign temp_13 = (((((((($signed(temp_9[1:0]) & temp_4) + temp_2[3:0]) ^ temp_11) ^ temp_2) | temp_10) * input_data) & (~input_data)) + temp_3[1:0]);
    assign temp_14 = temp_1 ? $signed((((($unsigned((($signed(temp_0) + temp_9) * temp_10[3:0])) + temp_0) * temp_10) ^ (~temp_8)) + (~temp_6))) : $signed(($unsigned(((((((($unsigned(input_data) - temp_4) | temp_8) | temp_4) ^ temp_10[15:0]) - temp_10) | temp_0) + temp_11)) | (~temp_13[1:0])));
    assign temp_15 = ((($signed((((temp_12 | temp_13) | (~temp_14)) | (~temp_12))) & temp_4) | temp_7) - temp_2);
    assign temp_16 = ($signed(($signed((temp_8 & temp_3)) + temp_4)) - (~temp_1));
    assign temp_17 = $signed(temp_13[14:0]);

    assign output_data = $signed(temp_10);

endmodule