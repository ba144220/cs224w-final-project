module top (
    input [3:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;

    assign temp_0 = (($signed(((($unsigned(($unsigned((input_data - input_data)) & input_data)) & input_data) ^ input_data) + input_data)) | input_data) - input_data);
    assign temp_1 = $signed(($unsigned(($unsigned(($signed(temp_0) ^ (~input_data))) * temp_0)) - input_data));
    assign temp_2 = ($signed(((($unsigned(($unsigned(($unsigned((temp_0[22:0] + input_data)) ^ temp_0)) * (~temp_1[8:0]))) | temp_1) & input_data) - input_data)) & input_data);
    assign temp_3 = temp_2;
    assign temp_4 = ((($signed((((temp_2 & temp_2) ^ input_data) + temp_2)) & temp_2) | temp_0) & input_data);
    assign temp_5 = $unsigned(((($unsigned((((temp_4 | temp_1) ^ temp_4) | temp_2)) | temp_4) + input_data) - temp_4));
    assign temp_6 = ($signed((($unsigned(((($unsigned(temp_3) | (~temp_2)) ^ temp_1) & temp_5)) * temp_1) | temp_3)) ^ temp_2);
    assign temp_7 = ((($unsigned((temp_1 + temp_0[12:0])) & temp_4) - temp_6) | temp_4);
    assign temp_8 = (((input_data * temp_0) + temp_3) - temp_0);
    assign temp_9 = ((((((($unsigned(temp_7) ^ temp_7) - temp_0) ^ temp_3[2:2]) * temp_0) + temp_3) + temp_1) & temp_6);
    assign temp_10 = $unsigned((((($unsigned(((temp_3 & temp_2) | temp_0)) - temp_7) | temp_8) | temp_2) - temp_3));
    assign temp_11 = temp_9 ? {2'b0, ((($signed((((temp_4 ^ temp_6) - temp_0) & temp_1)) | temp_3) & temp_7) + temp_7)} : ($signed(($signed(($unsigned(($unsigned(((temp_10 | temp_2) | temp_8)) * temp_0)) ^ temp_7)) ^ temp_1)) | temp_3);

    assign output_data = ((((((($signed(temp_1) & temp_9) * temp_10) & temp_10) - temp_7) - temp_3[2:2]) - temp_8) - temp_3[2:1]);

endmodule