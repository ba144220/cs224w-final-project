module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;

    assign temp_0 = $signed(input_data);
    assign temp_1 = ($unsigned((input_data - temp_0)) + input_data);
    assign temp_2 = ($signed((temp_1 | input_data)) & input_data);
    assign temp_3 = temp_2;
    assign temp_4 = $signed(input_data);
    assign temp_5 = ($signed(($unsigned((($signed(($signed(temp_0) & (~temp_2))) - temp_2) + temp_0)) | temp_1[25:17])) - temp_1);
    assign temp_6 = temp_1;
    assign temp_7 = input_data;
    assign temp_8 = ($signed((($signed(($unsigned(temp_7) & temp_4)) ^ temp_0) - temp_7)) + temp_2[29:0]);
    logic [21:0] expr_83560;
    assign expr_83560 = ($unsigned(temp_8) | temp_1[20:0]);
    assign temp_9 = expr_83560[3:0];
    assign temp_10 = $signed(($signed(($unsigned(($unsigned(($signed(temp_1[18:0]) & (~temp_4))) | (~temp_5))) - temp_7)) - temp_5));
    assign temp_11 = ($unsigned(($signed(($signed((temp_5 ^ temp_0)) | temp_8)) * input_data)) - (~temp_5));
    assign temp_12 = ($signed((temp_0 + temp_1[19:0])) + temp_1);
    logic [32:0] expr_968884;
    assign expr_968884 = ($unsigned((($unsigned(($unsigned(temp_5) ^ temp_7)) & temp_4) & temp_2)) * temp_4);
    assign temp_13 = expr_968884[11:0];
    assign temp_14 = ($unsigned(($unsigned(temp_9) | (~temp_3[2:0]))) | temp_10);
    assign temp_15 = (($unsigned(($unsigned(($unsigned(temp_2) | temp_1)) | temp_5[4:1])) * temp_1) * temp_7);

    logic [29:0] expr_819553;
    assign expr_819553 = ($unsigned((($unsigned(($unsigned(temp_11) & temp_1)) & temp_10[14:4]) ^ temp_1)) + temp_5);
    assign output_data = expr_819553[19:0];

endmodule