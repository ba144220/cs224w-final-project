module top (
    input [2:0] input_data,
    output [2:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;
    logic [17:0] temp_12;
    logic [2:0] temp_13;
    logic [1:0] temp_14;
    logic [23:0] temp_15;

    assign temp_0 = ((((($signed(input_data) | input_data) | input_data) & input_data) & input_data) | input_data);
    assign temp_1 = $unsigned(((((($unsigned(($signed((temp_0 * input_data)) * input_data)) ^ temp_0) + temp_0) | temp_0) ^ 24'd8371887) + temp_0[5:2]));
    assign temp_2 = temp_0;
    assign temp_3 = {17'b0, input_data};
    assign temp_4 = ($unsigned(input_data) > temp_1);
    assign temp_5 = ($unsigned(($signed((($signed(temp_1) + input_data) >= temp_2)) < temp_0[5:1])) & temp_3);
    assign temp_6 = temp_4;
    assign temp_7 = input_data[1:1] ? ($unsigned(($signed(($signed((temp_6[2:2] - input_data)) ^ temp_1)) ^ temp_6[2:2])) & input_data) : temp_5;
    assign temp_8 = (($unsigned(($signed((($signed(($signed((($unsigned(temp_6) * temp_2) | temp_1[6:0])) & input_data)) ^ input_data) & temp_3)) ^ (~temp_5))) | temp_2[10:5]) ^ temp_5);
    assign temp_9 = ((($unsigned(input_data) * temp_7) | temp_3[19:18]) ^ input_data);
    assign temp_10 = ((-24'd4072025 | temp_1) * temp_7[2:0]);
    assign temp_11 = ($signed(($signed((($unsigned(temp_2[8:0]) & input_data) * temp_6)) - temp_8)) * temp_6);
    assign temp_12 = ($signed(temp_3[19:4]) + temp_6);
    assign temp_13 = ($unsigned(($signed(temp_4[16:8]) & temp_10)) | temp_6);
    assign temp_14 = ($signed((($signed(((($signed(temp_12) | temp_10[10:0]) * temp_1) + temp_2)) & temp_5) - temp_3[19:5])) - temp_4[7:0]);
    assign temp_15 = temp_7;

    assign output_data = (($signed(((($unsigned(($signed(temp_15) - temp_15)) + temp_3) * temp_2) ^ temp_7)) >> (~temp_1)) + temp_1);

endmodule