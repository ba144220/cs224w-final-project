module top (
    input [3:0] input_data,
    output [2:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;
    logic [26:0] temp_10;
    logic [4:0] temp_11;
    logic [15:0] temp_12;
    logic [5:0] temp_13;
    logic [27:0] temp_14;
    logic [3:0] temp_15;
    logic [7:0] temp_16;
    logic [14:0] temp_17;
    logic [3:0] temp_18;

    assign temp_0 = (($unsigned((input_data | input_data)) == (~input_data)) + input_data);
    assign temp_1 = ($unsigned(($unsigned(input_data) | (~input_data))) & temp_0);
    assign temp_2 = ($unsigned((temp_0 ^ temp_1)) & input_data);
    assign temp_3 = ($unsigned(($signed((temp_1 - input_data)) ^ input_data)) + temp_2);
    assign temp_4 = (((($unsigned(input_data) & temp_0) + temp_0) | temp_1[3:2]) & (~temp_3));
    assign temp_5 = ($signed(input_data) | temp_0);
    assign temp_6 = ($signed(input_data) & (~input_data));
    assign temp_7 = ((input_data[3:1] + temp_1) | (~input_data[3:1]));
    assign temp_8 = ($signed(input_data) & temp_1);
    assign temp_9 = (($signed((temp_2[1:0] | input_data)) * temp_8) ^ temp_7);
    assign temp_10 = ((($unsigned((temp_0[25:5] > temp_1)) - input_data) <= temp_1) != temp_8);
    assign temp_11 = $signed(($unsigned(($unsigned((($signed(temp_6) + temp_6[11:0]) ^ temp_5)) + temp_7)) & temp_3[6:3]));
    assign temp_12 = temp_1;
    assign temp_13 = (($signed(($unsigned(input_data) ^ temp_4[23:0])) + (~temp_12)) + (~temp_8));
    assign temp_14 = ($signed((temp_4 > (~temp_2))) + temp_8);
    assign temp_15 = ($signed((($signed(temp_3) ^ (~temp_2)) ^ temp_6[13:7])) * temp_11);
    assign temp_16 = ($unsigned(temp_5[2:0]) - temp_6);
    assign temp_17 = ($unsigned(temp_4) >= temp_10);
    assign temp_18 = ($unsigned(((temp_16 + temp_7[2:2]) & (~temp_0))) + temp_16[7:5]);

    assign output_data = (temp_14 & (~temp_9));

endmodule