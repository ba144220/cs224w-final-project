module top (
    input [3:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;

    assign temp_0 = {17'b0, $signed(($unsigned((((input_data & input_data) & input_data) & input_data)) + (~input_data)))};
    assign temp_1 = $signed(($signed((($unsigned(($signed(temp_0) ^ temp_0)) - temp_0) | temp_0)) | input_data));
    assign temp_2 = $signed((($signed(($signed(temp_0) * temp_1)) & (~temp_0)) | temp_0));
    assign temp_3 = $signed(($signed(($signed(($unsigned((temp_1[8:0] - temp_2)) | temp_1)) & temp_1)) ^ (~temp_1)));
    assign temp_4 = temp_1;
    assign temp_5 = ($signed(($signed(temp_3) | temp_2)) * temp_2);
    assign temp_6 = ($unsigned(((temp_5 | (~temp_3)) - temp_5)) * temp_2);

    assign output_data = $unsigned(((($signed(temp_4) & temp_6) & temp_0) + temp_0));

endmodule