module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;

    assign temp_0 = input_data;
    assign temp_1 = ($unsigned((temp_0 * input_data)) ^ input_data);
    assign temp_2 = ($signed(($signed(($signed((($signed((($signed(temp_1) | input_data) ^ input_data)) * input_data) ^ input_data)) - input_data)) + input_data)) & input_data);
    assign temp_3 = 1'd0 ? ($signed((temp_0[5:3] - temp_1)) | input_data) : (($unsigned(($signed(($unsigned((((temp_1 * temp_2) ^ temp_0[5:4]) ^ input_data)) + temp_2)) + temp_1[23:3])) - temp_0) - input_data);
    assign temp_4 = (temp_0 * temp_3);
    assign temp_5 = (($signed(($unsigned(($unsigned(($unsigned(($unsigned(($signed(temp_0) ^ temp_3)) & input_data)) - temp_0)) & temp_2)) & input_data)) ^ temp_0) - input_data);
    assign temp_6 = (($unsigned(($unsigned((($unsigned((temp_3 - temp_3)) - temp_5) & temp_0)) + temp_3)) | temp_5[13:12]) ^ temp_5);
    assign temp_7 = temp_1 ? ($unsigned((($unsigned(temp_6) | temp_3[19:14]) ^ temp_6[2:2])) + temp_3) : (((($signed((temp_3 ^ temp_1)) * temp_0) * temp_1) * temp_5) + temp_1);
    assign temp_8 = (($unsigned(((((($signed(temp_1) & temp_3[19:15]) & input_data) * temp_1) - temp_2) ^ temp_5)) ^ temp_1) & temp_2);
    assign temp_9 = (($unsigned(((((temp_6 * temp_3[19:5]) * temp_4) + temp_5) - temp_4)) != temp_6[2:2]) >= temp_8);
    assign temp_10 = temp_1;
    assign temp_11 = temp_0 ? ($signed(((temp_1 & temp_7) | temp_0)) ^ temp_3) : (($unsigned((temp_6 | temp_10[23:5])) & temp_5) | temp_4);

    assign output_data = temp_3;

endmodule