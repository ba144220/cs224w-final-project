module top (
    input [3:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;

    assign temp_0 = ($unsigned(($unsigned(($unsigned(input_data) ^ input_data)) ^ input_data)) + input_data);
    logic [27:0] expr_695429;
    assign expr_695429 = ($signed(($unsigned(($unsigned(temp_0) & temp_0)) - input_data)) - temp_0);
    assign temp_1 = input_data[1:1] ? ($signed(($unsigned(input_data) | temp_0)) ^ input_data) : expr_695429[8:0];
    assign temp_2 = temp_1 ? ((($signed((($unsigned(($signed(($unsigned(temp_0) ^ temp_1)) | temp_0)) & input_data) - input_data)) & input_data) ^ temp_0) ^ input_data) : ($unsigned((($unsigned(input_data) & temp_0) <= temp_1)) ^ temp_1);
    assign temp_3 = $signed(($signed((($unsigned(($unsigned(($signed(input_data[2:0]) * temp_1)) * input_data[3:1])) * temp_0) - temp_0)) & input_data[2:0]));
    assign temp_4 = (input_data + input_data);
    assign temp_5 = (($unsigned(($unsigned(temp_4) | temp_1)) | temp_2) ^ temp_1);
    assign temp_6 = (($unsigned(temp_3) >> temp_3) ^ temp_5);
    assign temp_7 = ((temp_4 * temp_4) + temp_0[12:0]);
    assign temp_8 = input_data[0:0] ? (input_data | temp_1) : (temp_2 | temp_5);
    assign temp_9 = $signed(($unsigned(($signed(($unsigned(($unsigned((temp_7 * temp_4)) * temp_4)) ^ temp_2)) & temp_3)) + temp_4));
    assign temp_10 = ($unsigned(($unsigned(((($unsigned(temp_2) + temp_3) - temp_3) - temp_2[11:0])) ^ input_data)) + temp_7);
    assign temp_11 = temp_3 ? ((($unsigned(((($signed((temp_1 | temp_7)) & temp_8) ^ temp_3) * input_data)) + temp_6) & temp_0) - temp_0) : $signed(($signed(input_data) & temp_1[6:0]));
    assign temp_12 = $unsigned(temp_8);
    assign temp_13 = $signed(($signed(($signed(($signed(($unsigned((((temp_9 ^ temp_5) & temp_4) | temp_6)) ^ temp_7)) ^ temp_1)) | temp_3)) | temp_0));

    assign output_data = temp_13 ? $signed(($signed(($unsigned(($unsigned((($unsigned((temp_8 + temp_12)) + temp_11) - temp_3[2:2])) - temp_8)) & temp_0)) - temp_7)) : ((($unsigned(($unsigned((temp_0 + temp_0)) ^ temp_4)) | temp_7) - temp_3) ^ temp_8);

endmodule