module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;

    assign temp_0 = (($unsigned((($unsigned(input_data) * input_data) * input_data)) - input_data) | input_data);
    assign temp_1 = ($unsigned((($unsigned(($unsigned(((input_data + temp_0) * temp_0[2:0])) - temp_0)) * input_data) + temp_0)) + temp_0);
    assign temp_2 = (($signed(($signed(((($signed((input_data * temp_0)) & input_data) | input_data) * input_data)) - temp_0)) & input_data) - temp_1);
    assign temp_3 = $unsigned((($unsigned(($unsigned(((((($unsigned(($signed(($signed(temp_1[7:0]) | input_data)) * input_data)) * input_data) * input_data) & input_data) - temp_1[25:0]) | temp_0)) & input_data)) * input_data) * input_data));
    assign temp_4 = ((($unsigned((($unsigned(((($unsigned((($signed(($signed(((temp_2 ^ input_data) & temp_1)) * temp_0[6:3])) | temp_0) ^ temp_0)) | temp_3) ^ temp_3[3:0]) * input_data)) + temp_1) | input_data)) - temp_3) - input_data) * input_data);
    logic [39:0] expr_827813;
    assign expr_827813 = ($signed(($unsigned(((($signed((($signed((($unsigned((input_data[5:1] * temp_4[2:0])) | temp_2) ^ input_data[5:1])) & temp_3) + temp_4)) | temp_0) ^ temp_1) ^ temp_2)) - temp_2)) & temp_2);
    assign temp_5 = expr_827813[4:0];
    assign temp_6 = ($unsigned((temp_1 != temp_3)) < temp_1);
    assign temp_7 = ($signed(((($signed(((($unsigned(((temp_4 * input_data) - input_data)) * input_data) - temp_5[2:0]) | input_data)) + input_data) ^ input_data) & temp_3)) | temp_6);
    logic [33:0] expr_56046;
    assign expr_56046 = (((($unsigned(($unsigned((temp_3 + temp_4)) - temp_3)) ^ temp_7) * temp_2) ^ temp_2) ^ input_data);
    assign temp_8 = expr_56046[18:0];
    assign temp_9 = (($signed(((($unsigned((($signed(($unsigned(($signed((temp_4 & temp_3)) * temp_6)) - temp_3)) - temp_5) ^ temp_8[18:10])) - temp_6) ^ temp_6) + temp_8[8:0])) ^ temp_6) * temp_5);
    assign temp_10 = (($unsigned((((temp_8 - temp_1[21:0]) - temp_2) + temp_0)) + temp_4) - temp_6[1:0]);
    assign temp_11 = (temp_3 - temp_1[25:1]);
    assign temp_12 = (($signed(($signed(((temp_8[2:0] + temp_2) ^ temp_9)) + temp_4)) | temp_7) | temp_8);
    assign temp_13 = (($signed(($unsigned(($unsigned(($signed(temp_5) >= temp_5)) == temp_2)) + temp_10)) & temp_11) < temp_2);

    assign output_data = temp_6;

endmodule