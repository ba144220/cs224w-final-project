module top (
    input [2:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;
    logic [1:0] temp_17;
    logic [16:0] temp_18;

    assign temp_0 = {3'b0, $signed((input_data + input_data))};
    assign temp_1 = ((input_data < temp_0) + temp_0);
    assign temp_2 = $signed((((temp_0 * input_data) - (~temp_0)) * input_data));
    assign temp_3 = $signed((((10'd909 * temp_1) & temp_1) - temp_0));
    assign temp_4 = input_data;
    assign temp_5 = {2'b0, input_data};
    assign temp_6 = (temp_2 * temp_4);
    assign temp_7 = (26'd63247293 ^ temp_3);
    assign temp_8 = ((temp_2 + input_data) & temp_0);
    assign temp_9 = ($unsigned(temp_5) & input_data);
    assign temp_10 = ((input_data - temp_8) > input_data);
    assign temp_11 = (((temp_4 - 24'd5917355) ^ temp_0[6:3]) != temp_8);
    assign temp_12 = input_data;
    assign temp_13 = $signed((((temp_10 | temp_12) * temp_1) * temp_4));
    assign temp_14 = (temp_1 + temp_7);
    assign temp_15 = (temp_3 | input_data);
    assign temp_16 = $unsigned(((temp_11 + temp_2) * temp_8));
    assign temp_17 = temp_8;
    assign temp_18 = $signed(temp_9);

    assign output_data = temp_17;

endmodule