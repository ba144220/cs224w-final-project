module top (
    input [2:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;
    logic [25:0] temp_16;

    assign temp_0 = input_data[0:0] ? (($signed((((((($unsigned((($signed((input_data ^ 25'd4233809)) + input_data) | input_data)) + input_data) | input_data) & 25'd6550931) * input_data) - (~input_data)) | input_data)) * input_data) ^ (~input_data)) : input_data;
    assign temp_1 = (($signed(((($unsigned(($unsigned((((temp_0 + temp_0) - (~input_data)) + input_data)) * temp_0)) | temp_0) & input_data) - input_data)) & (~input_data)) ^ temp_0);
    assign temp_2 = ((($unsigned((((((($signed(temp_0[20:0]) * input_data) ^ temp_1) * temp_0) * temp_1) ^ temp_1) + temp_0)) | input_data) ^ temp_1) - input_data);
    assign temp_3 = ($unsigned(((($unsigned(($unsigned((($signed(((3'd4 + (~temp_1)) | (~temp_2))) - temp_1) - temp_1)) | (~temp_0))) | (~temp_1)) ^ temp_0) & temp_2)) * temp_0);
    assign temp_4 = ((((((((($unsigned(temp_3) | temp_2) | temp_2) & temp_0[24:12]) & temp_1[8:3]) & temp_0) * input_data) - temp_3) * input_data) ^ temp_0);
    assign temp_5 = temp_2;
    assign temp_6 = ($unsigned(temp_4) ^ temp_3);
    assign temp_7 = temp_5 ? (($signed(($unsigned(($unsigned(($signed(((($unsigned(((temp_0[15:0] ^ input_data) ^ temp_2[12:4])) & temp_6[11:0]) ^ input_data) - temp_6)) ^ temp_3)) ^ temp_0)) & temp_5)) & temp_6) | temp_3) : (((((temp_1 - temp_1) - temp_5) * temp_3) + (~temp_4)) + input_data);
    assign temp_8 = (temp_0 + temp_5);
    assign temp_9 = ($signed(((($signed((($unsigned(((((temp_7 | input_data[1:0]) & input_data[1:0]) | temp_2) | temp_8)) * temp_0) ^ input_data[2:1])) | temp_1) - temp_5) + temp_4)) & temp_4);
    assign temp_10 = temp_7 ? ($signed((($unsigned((((($signed(($unsigned((((temp_6 ^ temp_7) - temp_8[11:0]) - temp_8)) & input_data)) - temp_8) & temp_7) | temp_0) ^ temp_5)) + temp_0) * temp_8)) - temp_4) : ($unsigned(((input_data | (~temp_4)) + temp_4)) - temp_8);
    logic [33:0] expr_702472;
    assign expr_702472 = ($unsigned((($unsigned(((((($unsigned(((input_data + temp_9[1:1]) * temp_9)) ^ (~temp_3)) * temp_8) - temp_4) & temp_1) | temp_10)) - temp_8) + temp_3)) & temp_9);
    assign temp_11 = expr_702472[31:0];
    assign temp_12 = ((($signed(($signed((($unsigned((((temp_2 - temp_1) ^ temp_9) * temp_11)) + temp_10) * temp_10)) | temp_4)) + (~temp_3)) + temp_3) | temp_2);
    assign temp_13 = ($signed(($signed(($signed((((((temp_4 + temp_7) | temp_11) << temp_5) << temp_5) - (~temp_10))) + temp_3)) | temp_9)) | temp_11);
    assign temp_14 = (temp_13 ^ (~temp_6));
    assign temp_15 = ($unsigned(($signed(temp_1) - temp_6)) & temp_2);
    assign temp_16 = ((($unsigned(((temp_5 * temp_4) & temp_13[24:9])) != (~temp_5)) * temp_6) ^ temp_13);

    assign output_data = (($unsigned(($signed((($signed(temp_3) * temp_10) * (~temp_2[6:0]))) + temp_11)) * temp_11) & temp_15);

endmodule