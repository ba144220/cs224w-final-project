module top (
    input [4:0] input_data,
    output [9:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;
    logic [0:0] temp_13;
    logic [28:0] temp_14;
    logic [17:0] temp_15;

    assign temp_0 = (((input_data + input_data) & input_data) >> input_data);
    assign temp_1 = input_data[0:0] ? ((temp_0 | input_data) & input_data) : (((((input_data ^ (~temp_0)) + (~temp_0)) - temp_0) * input_data) ^ (~temp_0));
    assign temp_2 = ((((((((temp_0 | temp_0) + input_data) + temp_0) | temp_1[6:0]) ^ (~temp_1)) & temp_0) | temp_0) & input_data);
    assign temp_3 = {24'b0, $signed(temp_2)};
    assign temp_4 = temp_2 ? ((((input_data | temp_0) & temp_3) * temp_3[31:7]) | input_data) : (((((((((((((input_data + temp_1) * temp_2) ^ input_data) & input_data) & temp_1) | (~input_data)) * temp_0[1:0]) - temp_3) + temp_3) ^ temp_0) * (~input_data)) * input_data) | input_data);
    assign temp_5 = temp_3[19:0] ? ((((((((((31'd1300556176 - temp_4) - (~temp_2[7:1])) * temp_1) ^ temp_1) | input_data) ^ temp_2) ^ input_data) ^ input_data) & temp_4) - (~temp_0)) : (((((((((input_data - temp_1) & input_data) & input_data) ^ temp_1[3:0]) * temp_1) ^ temp_3) | temp_1) + temp_3) ^ input_data);
    assign temp_6 = ((input_data & input_data) & temp_2);
    assign temp_7 = ((((((((((temp_0 | temp_5) - temp_2) - temp_3) - temp_0[4:1]) ^ input_data) | temp_6[24:15]) | temp_6) & temp_0) ^ temp_3) * (~temp_3));
    assign temp_8 = $unsigned((((((((((((((temp_1 ^ input_data) ^ temp_6) | temp_4) & input_data) + (~temp_6[3:0])) | temp_2) - temp_3) | temp_7) ^ input_data) | temp_7) | temp_0) - temp_3[24:0]) & temp_2));
    assign temp_9 = (((temp_1 & input_data) - temp_7) * temp_4);
    assign temp_10 = (((temp_6 * temp_1) & temp_6) ^ temp_0[2:0]);
    assign temp_11 = temp_4[28:2] ? ((((((((temp_1 >> temp_4) | input_data) * temp_9) << temp_8) - temp_1) + (~temp_8)) + temp_2) | (~temp_5[2:0])) : ((((temp_4[27:0] - temp_3) | temp_2) | temp_8[3:0]) & temp_1);
    assign temp_12 = (((((temp_8[1:0] - temp_11) & temp_5) | temp_2[4:0]) - temp_11) * temp_5);
    assign temp_13 = ((((((temp_8 - temp_10) - temp_2) & temp_4) - temp_10) + temp_4[28:18]) & (~temp_9));
    assign temp_14 = ((((temp_13 ^ temp_12) | temp_8) | temp_2) & temp_9[14:0]);
    assign temp_15 = (temp_12 & temp_6[24:12]);

    assign output_data = ((temp_13 ^ temp_13) ^ (~temp_15));

endmodule