module top (
    input [6:0] input_data,
    output [11:0] output_data
);

    logic [1:0] temp_0;
    logic [29:0] temp_1;
    logic [15:0] temp_2;
    logic [3:0] temp_3;
    logic [10:0] temp_4;
    logic [7:0] temp_5;
    logic [23:0] temp_6;
    logic [30:0] temp_7;
    logic [15:0] temp_8;
    logic [24:0] temp_9;
    logic [6:0] temp_10;
    logic [15:0] temp_11;
    logic [0:0] temp_12;
    logic [13:0] temp_13;
    logic [26:0] temp_14;
    logic [17:0] temp_15;
    logic [11:0] temp_16;
    logic [24:0] temp_17;

    assign temp_0 = $signed(-2'd1);
    assign temp_1 = {22'b0, $signed((input_data - input_data))};
    assign temp_2 = ((($unsigned((16'd40116 & (~input_data))) + input_data) | input_data) + input_data);
    assign temp_3 = $unsigned(((($unsigned(((temp_1[29:11] | input_data[5:2]) + temp_1)) * input_data[3:0]) + (~temp_2)) ^ temp_1));
    assign temp_4 = ((temp_3 - input_data) * temp_3[3:3]);
    assign temp_5 = ((temp_0 ^ temp_0) & temp_2);
    assign temp_6 = ((temp_2 ^ input_data) * input_data);
    assign temp_7 = temp_3 ? ((((temp_4 ^ (~input_data)) ^ (~temp_5)) - temp_1) ^ temp_4) : $unsigned(input_data);
    logic [25:0] expr_660032;
    assign expr_660032 = ((input_data & temp_6) * input_data);
    assign temp_8 = expr_660032[15:0];
    assign temp_9 = $unsigned(((((temp_4 & input_data) * (~temp_5)) + (~temp_7[30:5])) | temp_3));
    assign temp_10 = (((input_data - (~temp_8)) * temp_9[24:18]) ^ temp_0);
    assign temp_11 = ($signed(((temp_4 * input_data) & input_data)) * temp_6);
    logic [30:0] expr_95879;
    assign expr_95879 = (temp_9 ^ temp_1);
    assign temp_12 = temp_1 ? temp_1[29:10] : expr_95879[0:0];
    logic [30:0] expr_556481;
    assign expr_556481 = ((((temp_0 | temp_8) + temp_4) * (~temp_6)) ^ temp_1);
    assign temp_13 = expr_556481[13:0];
    assign temp_14 = temp_0 ? $signed((((temp_10 ^ temp_5) & temp_11) * (~temp_9))) : $signed(((($signed(temp_0) | (~input_data)) * temp_13[13:5]) * (~temp_0[1:1])));
    assign temp_15 = (((((temp_2 | temp_1) - temp_4) - (~temp_0)) + temp_10[6:5]) | (~temp_1));
    assign temp_16 = (((temp_13 + temp_6) - (~temp_3)) & temp_14);
    assign temp_17 = ((temp_3 * temp_10) & temp_7);

    assign output_data = temp_17[10:0];

endmodule