module top (
    input [2:0] input_data,
    output [4:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;
    logic [1:0] temp_17;

    assign temp_0 = ($unsigned((input_data + input_data)) - input_data);
    assign temp_1 = ($signed(($signed(((input_data | temp_0) + temp_0)) ^ temp_0)) | temp_0);
    assign temp_2 = (temp_0 ^ temp_1);
    logic [26:0] expr_772927;
    assign expr_772927 = ($signed(temp_2[2:0]) & temp_1);
    assign temp_3 = input_data[1:1] ? expr_772927[9:0] : (input_data * 10'd838);
    assign temp_4 = (input_data - temp_2);
    assign temp_5 = ($signed(($signed(temp_0[6:2]) | input_data)) * input_data);
    assign temp_6 = ($unsigned(temp_2[30:6]) != temp_4);
    assign temp_7 = ($unsigned(((input_data - temp_2) & temp_0)) - temp_0);
    assign temp_8 = ((input_data + input_data) ^ 19'd205366);
    assign temp_9 = (($unsigned(temp_7) + temp_0) - temp_6);
    assign temp_10 = ((temp_9 & temp_7) * temp_1);
    assign temp_11 = ((($unsigned((temp_2 * temp_0)) ^ temp_1) - temp_7) | input_data);
    assign temp_12 = ($signed(((($unsigned(temp_6) & temp_0) & input_data) ^ input_data)) & temp_7);
    assign temp_13 = (($signed(((temp_8 - temp_5) | input_data)) ^ temp_8[18:18]) * temp_1);
    assign temp_14 = ($unsigned(temp_10[13:0]) - temp_1);
    assign temp_15 = (((temp_3 ^ temp_10) & temp_13) ^ temp_1);
    assign temp_16 = ($unsigned((temp_7 ^ temp_4)) + temp_7);
    assign temp_17 = ((temp_12 + temp_16) & temp_6[1:0]);

    assign output_data = (($signed((temp_8[18:13] * temp_9)) - temp_2) + temp_10[10:0]);

endmodule