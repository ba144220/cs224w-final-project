module top (
    input [5:0] input_data,
    output [39:0] output_data
);

    logic [23:0] temp_0;
    logic [17:0] temp_1;
    logic [8:0] temp_2;
    logic [11:0] temp_3;
    logic [0:0] temp_4;
    logic [21:0] temp_5;
    logic [29:0] temp_6;
    logic [5:0] temp_7;
    logic [21:0] temp_8;
    logic [2:0] temp_9;
    logic [24:0] temp_10;
    logic [10:0] temp_11;
    logic [28:0] temp_12;
    logic [27:0] temp_13;
    logic [10:0] temp_14;
    logic [10:0] temp_15;
    logic [15:0] temp_16;
    logic [3:0] temp_17;

    assign temp_0 = ((((input_data ^ input_data) & input_data) * (~input_data)) & input_data);
    assign temp_1 = ((((temp_0 * temp_0) - temp_0) + temp_0) != temp_0);
    assign temp_2 = ($signed((($unsigned(((($signed(temp_1) | input_data) * temp_0) & input_data)) | input_data) | temp_1)) - temp_0);
    assign temp_3 = ((temp_0 + temp_1) - temp_1);
    assign temp_4 = (($unsigned((((input_data[1:1] - temp_3) + 1'd1) | temp_0)) - temp_0) ^ temp_2);
    assign temp_5 = ($signed((($unsigned((temp_3 + temp_1[17:16])) ^ input_data) & input_data)) & input_data);
    assign temp_6 = {25'b0, temp_5[21:17]};
    assign temp_7 = (($signed(((input_data > input_data) * temp_6)) + input_data) ^ temp_2);
    assign temp_8 = (((temp_5 + temp_5) & input_data) * temp_6);
    assign temp_9 = ((temp_5[5:0] * temp_1) & input_data[3:1]);
    assign temp_10 = ((((input_data * temp_0) + temp_2) - temp_5) | temp_1);
    assign temp_11 = ((((input_data & temp_5) - temp_2) & input_data) ^ temp_2[4:0]);
    assign temp_12 = temp_11[3:0];
    assign temp_13 = ((($signed(((temp_12 - temp_0) - temp_10)) * temp_12) | temp_1[17:15]) * temp_2);
    assign temp_14 = ((((($unsigned(temp_0) != temp_5) * temp_9) & temp_5) <= temp_7) - temp_5);
    assign temp_15 = (((temp_1 & temp_4) & temp_0) + temp_9);
    assign temp_16 = ((temp_6 ^ temp_10) | temp_15);
    assign temp_17 = ((((temp_13 | temp_9) * temp_5) | temp_11) ^ temp_15);

    assign output_data = temp_2;

endmodule