module top (
    input [2:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;
    logic [25:0] temp_16;
    logic [5:0] temp_17;
    logic [31:0] temp_18;

    assign temp_0 = input_data;
    assign temp_1 = $unsigned((temp_0 & input_data));
    assign temp_2 = $unsigned((($signed(($signed(((((((temp_1 - input_data) & input_data) ^ temp_0) + temp_1) + (~temp_0)) & temp_0)) & temp_0)) * temp_1) & input_data));
    assign temp_3 = $unsigned(input_data);
    assign temp_4 = (input_data + temp_3);
    assign temp_5 = (((((((temp_0[24:20] | input_data) ^ input_data) & input_data) + input_data) | temp_2) * input_data) | input_data);
    assign temp_6 = (((((temp_3 | input_data) & input_data) | temp_5) ^ temp_1) + input_data);
    assign temp_7 = (((($unsigned(((((($unsigned(temp_3) | temp_4) + input_data) - input_data) * temp_0) & temp_5)) - temp_1[1:0]) - temp_2) ^ input_data) - temp_6);
    assign temp_8 = (((((temp_5 - temp_7) | temp_4) & temp_1) * temp_0) - temp_2);
    assign temp_9 = $signed((((((((((input_data[2:1] ^ temp_2) & temp_0) + temp_3) - temp_0) * temp_7) * temp_1) & temp_8) + temp_4) - (~2'd1)));
    assign temp_10 = ($unsigned(($signed(((temp_1 + input_data) ^ input_data)) - temp_5)) + temp_7);
    assign temp_11 = input_data[2:2] ? (((temp_7 - temp_1) & input_data) & temp_8) : ((((((((($signed(temp_4[3:0]) | temp_3) * temp_6) + (~temp_8)) + input_data) | temp_2[8:0]) - temp_1[6:0]) & temp_7) + temp_7) ^ temp_8);
    assign temp_12 = $signed((((((((((input_data | temp_8) * temp_0) | input_data) - temp_1) + temp_2) & temp_6[6:0]) & temp_9[1:0]) + temp_7) * temp_7));
    assign temp_13 = ((temp_3 ^ (~input_data)) * input_data);
    assign temp_14 = (((temp_2 * temp_7) | input_data) & temp_0);
    assign temp_15 = (((($unsigned(temp_10) & input_data) - temp_5) + temp_13) ^ -13'd3127);
    assign temp_16 = $signed((((((temp_10 ^ (~temp_9)) + temp_9) - temp_4) ^ temp_4) | temp_10));
    assign temp_17 = $unsigned(temp_16[25:1]);
    assign temp_18 = (((((temp_17 & temp_12) & temp_3) | temp_1) - temp_12) + temp_7);

    assign output_data = $unsigned(((temp_5 + temp_12) ^ temp_8));

endmodule