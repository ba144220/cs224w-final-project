module top (
    input [3:0] input_data,
    output [3:0] output_data
);

    logic [16:0] temp_0;
    logic [2:0] temp_1;
    logic [0:0] temp_2;
    logic [9:0] temp_3;
    logic [30:0] temp_4;
    logic [23:0] temp_5;
    logic [20:0] temp_6;
    logic [1:0] temp_7;
    logic [17:0] temp_8;
    logic [31:0] temp_9;
    logic [12:0] temp_10;
    logic [26:0] temp_11;

    assign temp_0 = ($signed(($signed(($unsigned(($signed((($signed(((input_data ^ input_data) + input_data)) + input_data) ^ input_data)) | input_data)) * input_data)) | input_data)) | input_data);
    assign temp_1 = ($unsigned(($unsigned(($signed(($unsigned(($unsigned(temp_0) ^ input_data[3:1])) ^ input_data[3:1])) ^ input_data[2:0])) - temp_0)) | temp_0);
    assign temp_2 = ($signed(($unsigned(($signed(($signed(($unsigned(($signed((($signed(($unsigned(($signed(input_data[3:3]) ^ temp_1)) | temp_1)) * (~temp_1[2:1])) | temp_1)) - temp_0)) ^ input_data[1:1])) ^ input_data[3:3])) - input_data[3:3])) + (~input_data[2:2]))) * temp_1);
    assign temp_3 = ($unsigned(($signed(input_data) << temp_0)) - temp_1[2:1]);
    assign temp_4 = ($signed(($unsigned(($unsigned(($unsigned((($signed(($signed(($signed(($signed((($signed(temp_1) | temp_3) | temp_1)) ^ (~temp_1))) + temp_0)) | temp_2)) & temp_0) ^ temp_2)) | input_data)) ^ input_data)) ^ temp_0)) * temp_0);
    assign temp_5 = ($unsigned((($unsigned(((($unsigned(((temp_4 & input_data) & temp_1)) + temp_3) & temp_3) * temp_2)) + input_data) + temp_3)) + temp_3);
    logic [27:0] expr_978979;
    assign expr_978979 = $unsigned(($unsigned((($signed(($signed(temp_5) - temp_0)) & (~temp_1[2:2])) * temp_1)) - temp_0));
    assign temp_6 = expr_978979[20:0];
    assign temp_7 = (temp_6 & temp_6[18:0]);
    assign temp_8 = ($signed(($unsigned(temp_1) | input_data)) * temp_4);
    assign temp_9 = temp_7 ? temp_3[9:5] : ($unsigned(($signed((temp_5 & input_data)) + temp_1[2:1])) + temp_8);
    assign temp_10 = (($signed(($unsigned(($signed(($signed(($unsigned(($signed(($signed(temp_0) ^ (~input_data))) ^ temp_0)) ^ temp_1)) + temp_8)) ^ temp_1)) - temp_4)) | temp_6) & temp_2);
    assign temp_11 = (($unsigned(($signed(($signed(temp_3) & temp_1[2:2])) & temp_5)) - temp_9) & (~temp_7[1:1]));

    assign output_data = $unsigned(($signed((($signed(($unsigned(($unsigned((($signed(($signed(($signed(($signed(temp_11) ^ temp_5)) + temp_5)) | temp_6)) ^ (~temp_0[7:0])) - temp_8)) ^ temp_2)) ^ temp_7)) & temp_11) + temp_10)) - temp_11));

endmodule