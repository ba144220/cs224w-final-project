module top (
    input [2:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;

    assign temp_0 = (((25'd27357858 > input_data) - input_data) - (~input_data));
    assign temp_1 = (temp_0 & input_data);
    assign temp_2 = ((((input_data * temp_1) ^ input_data) + temp_1) + (~temp_0));
    logic [24:0] expr_911111;
    assign expr_911111 = ($unsigned(($unsigned(($unsigned(input_data) - temp_0[22:0])) >> input_data)) - input_data);
    assign temp_3 = expr_911111[2:0];
    assign temp_4 = (($signed((($unsigned(temp_0) & input_data) - input_data)) & (~input_data)) ^ temp_0);
    assign temp_5 = (($signed(((temp_4[5:5] * input_data) | temp_2)) * input_data) * temp_3);
    assign temp_6 = ((input_data * (~temp_3)) * input_data);
    assign temp_7 = $signed(((($signed((input_data * temp_0)) & input_data) + (~temp_6)) * input_data));
    assign temp_8 = temp_5;
    assign temp_9 = (((((temp_6 + temp_3) + temp_2) ^ temp_1) - (~temp_3)) & temp_4);
    assign temp_10 = {2'b0, (((temp_2 & input_data) | temp_8) & temp_1[8:6])};
    assign temp_11 = (((((temp_2 >= temp_1) ^ input_data) * temp_7) ^ temp_10[5:0]) == temp_0);
    assign temp_12 = temp_4;
    assign temp_13 = temp_9;
    assign temp_14 = $unsigned((((($signed(temp_2) + temp_12) - temp_0[23:0]) + input_data) + temp_3));
    assign temp_15 = (($signed((temp_6 - temp_10)) | (~temp_0)) & temp_2);

    assign output_data = (temp_6 ^ temp_15);

endmodule