module top (
    input [5:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;

    assign temp_0 = input_data;
    assign temp_1 = $unsigned(temp_0);
    assign temp_2 = ($signed(input_data) | input_data);
    assign temp_3 = $signed(($signed(($signed(($unsigned(($signed(temp_0[24:23]) * temp_2)) | temp_2)) - temp_1)) + temp_2[12:3]));
    logic [27:0] expr_629823;
    assign expr_629823 = $signed(($signed(($signed(($unsigned(($unsigned(($signed(($signed(temp_0[24:3]) ^ temp_2)) - temp_1)) * temp_3)) | temp_2)) & temp_3)) ^ (~temp_3)));
    assign temp_4 = expr_629823[5:0];
    assign temp_5 = $signed(temp_4);
    assign temp_6 = (($unsigned((temp_5 < temp_2[7:0])) != temp_4) - temp_2);
    assign temp_7 = ($signed(($unsigned(($unsigned(($unsigned(((($unsigned(($unsigned(temp_4) - temp_4[5:2])) & temp_4) * temp_5) ^ temp_1)) + temp_3[1:0])) - temp_1[8:8])) | temp_4)) + (~temp_5));

    assign output_data = ($signed(($signed(($signed(($unsigned(($signed(temp_5) < temp_2)) * temp_5)) * temp_5)) - temp_2)) > temp_0);

endmodule