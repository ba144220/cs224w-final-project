module top (
    input [3:0] input_data,
    output [9:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;
    logic [26:0] temp_10;
    logic [4:0] temp_11;
    logic [15:0] temp_12;
    logic [5:0] temp_13;
    logic [27:0] temp_14;
    logic [3:0] temp_15;
    logic [7:0] temp_16;
    logic [14:0] temp_17;

    assign temp_0 = {22'b0, input_data};
    assign temp_1 = $unsigned(((((((((input_data * temp_0) * temp_0) + input_data) + temp_0) ^ temp_0) + (~input_data)) ^ input_data) ^ temp_0));
    assign temp_2 = $signed((((((((input_data | temp_1) + temp_0) * (~temp_1)) | input_data) ^ input_data) & temp_0) + (~temp_0)));
    assign temp_3 = (((((temp_1 - temp_1) - input_data) | temp_2) - temp_0) - input_data);
    assign temp_4 = (((((((input_data * temp_0) | (~input_data)) ^ temp_3) ^ temp_3) - temp_3) ^ input_data) ^ input_data);
    logic [27:0] expr_102493;
    assign expr_102493 = $signed(((((temp_4 ^ temp_3) | temp_1) + input_data) | temp_4));
    assign temp_5 = expr_102493[3:0];
    assign temp_6 = ((((((((temp_2 <= temp_2) != temp_2) < temp_3) | input_data) ^ temp_1) > temp_5) ^ temp_2) > (~input_data));
    assign temp_7 = (input_data[2:0] & input_data[3:1]);
    logic [16:0] expr_768690;
    assign expr_768690 = $signed(((((temp_1 + (~6'd8)) + temp_6) - input_data) * temp_3));
    assign temp_8 = expr_768690[5:0];
    assign temp_9 = (((temp_6 & input_data) ^ (~temp_2)) + temp_4);
    assign temp_10 = ((((temp_0 | (~temp_0)) & (~temp_4)) * input_data) ^ temp_9);
    assign temp_11 = (((((((temp_0 | temp_8[5:0]) + (~input_data)) ^ (~temp_1)) | temp_7) | (~temp_8[4:0])) * temp_3) + temp_10);
    assign temp_12 = ((((temp_7 ^ temp_7) + input_data) + temp_1) - input_data);
    assign temp_13 = $signed(((((((((temp_7 + temp_7) & (~temp_5[2:0])) - temp_11) | (~temp_6)) ^ temp_2) * temp_6) | temp_11[4:0]) ^ temp_7[1:0]));
    assign temp_14 = $signed(((((((temp_6[11:0] - temp_8) & (~temp_8)) - temp_12) & temp_3) * (~temp_8)) - temp_10));
    assign temp_15 = $signed((((((((temp_14 & input_data) ^ temp_13) | temp_0) * (~input_data)) + (~temp_9)) | temp_7) | temp_3[4:0]));
    assign temp_16 = $unsigned(((((temp_15[2:0] ^ temp_12) - temp_6) * temp_15) + temp_4));
    assign temp_17 = $signed((((((temp_10 | temp_1) & temp_0[3:0]) + temp_6) + temp_15) ^ temp_0));

    assign output_data = temp_6 ? (((((temp_1 * temp_8) + temp_0) & temp_8) + temp_9) * temp_14) : (temp_17 + temp_2);

endmodule