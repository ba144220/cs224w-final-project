module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;

    assign temp_0 = ($signed(input_data) ^ input_data);
    assign temp_1 = ($signed(($signed(input_data) - input_data)) * input_data);
    assign temp_2 = {5'b0, temp_1};
    assign temp_3 = ($signed(($signed(($unsigned(($unsigned(($signed(temp_2) - input_data)) - temp_0[6:3])) ^ input_data)) & input_data)) - temp_2);
    assign temp_4 = $signed(input_data);
    assign temp_5 = ($signed(temp_2) | temp_3);
    assign temp_6 = ($signed(($signed((temp_2 - temp_2[2:0])) + input_data[1:0])) | input_data[3:2]);
    assign temp_7 = ($unsigned(($unsigned(($unsigned((($signed(temp_3[5:0]) ^ temp_0) - temp_3)) + temp_1[9:0])) - temp_1[20:0])) & input_data);
    assign temp_8 = ($unsigned(($signed(input_data) + temp_7)) & temp_1);
    assign temp_9 = ($unsigned(temp_1) - (~temp_2));
    assign temp_10 = temp_1;
    assign temp_11 = (($unsigned(($unsigned(($unsigned(($signed(temp_8) >= temp_8)) ^ temp_5[1:0])) | temp_5)) == temp_2) <= temp_1);

    assign output_data = temp_1;

endmodule