module top (
    input [4:0] input_data,
    output [36:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;

    assign temp_0 = ($unsigned(($unsigned(($unsigned(((($signed((($signed(((((input_data & input_data) - (~input_data)) + input_data) - input_data)) & input_data) * input_data)) ^ input_data) ^ input_data) - input_data)) | input_data)) - (~input_data))) - input_data);
    assign temp_1 = ($signed((($signed(($unsigned((((((temp_0 | temp_0) | temp_0) | (~input_data)) * temp_0) + temp_0[4:2])) - (~input_data))) + temp_0[4:2]) | input_data)) & temp_0);
    assign temp_2 = ($unsigned(($signed(($signed(($signed((($signed(($unsigned(((((($unsigned((temp_0 ^ temp_1)) | (~temp_0)) * temp_0) * temp_1) | temp_1) | temp_0)) - temp_1)) + temp_1) + input_data)) | temp_0[1:0])) - temp_1)) | temp_1[4:0])) - temp_1[13:0]);
    assign temp_3 = ($signed(($unsigned(((((((temp_0[4:1] + temp_0) & temp_0[1:0]) | input_data) - temp_0[3:0]) & temp_0[3:0]) + temp_2)) * (~temp_2))) & temp_2);
    assign temp_4 = {11'b0, ($unsigned(($unsigned(($unsigned(($unsigned(temp_0[4:2]) << temp_0[4:1])) * temp_2[6:0])) ^ (~temp_2[2:0]))) ^ temp_1)};
    assign temp_5 = $signed(((((($signed(((($unsigned((($unsigned(($unsigned((temp_4 * temp_3[21:0])) + temp_2)) | temp_4[16:0]) ^ temp_1)) & (~temp_4)) + temp_2[7:0]) * temp_4)) + temp_4) + temp_3) ^ temp_4) + temp_1) + temp_1));

    assign output_data = (((temp_3 * temp_1) | temp_0[2:0]) * temp_1);

endmodule