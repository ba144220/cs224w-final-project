module top (
    input [3:0] input_data,
    output [9:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;
    logic [1:0] temp_17;
    logic [16:0] temp_18;

    assign temp_0 = $signed((input_data - input_data));
    assign temp_1 = ($signed(((((($signed(temp_0) | temp_0) + temp_0) * temp_0[2:0]) - temp_0) ^ (~temp_0))) * temp_0);
    assign temp_2 = ($unsigned(($signed(((temp_1 | input_data) * input_data)) - temp_0[1:0])) - temp_1);
    assign temp_3 = ($signed(temp_1) & input_data);
    assign temp_4 = ((temp_3 != temp_3) * temp_3);
    assign temp_5 = ($unsigned(((input_data + temp_4) - temp_3)) + temp_1[9:0]);
    assign temp_6 = {1'b0, ($unsigned(input_data[2:1]) <= temp_0[5:0])};
    assign temp_7 = input_data[2:2] ? (((((($signed(input_data) * temp_6) * temp_3) - temp_6[1:1]) ^ (~temp_3)) - temp_2[30:26]) + temp_3) : ($unsigned((((input_data | temp_4) ^ temp_3[3:0]) * input_data)) + temp_1);
    assign temp_8 = temp_1 ? (((temp_1 ^ temp_4) & temp_4) & input_data) : ((temp_5 + temp_1) * input_data);
    assign temp_9 = {3'b0, $signed(($signed(temp_6) <= (~temp_8)))};
    assign temp_10 = (($signed(temp_2) ^ temp_8[18:18]) * temp_1);
    assign temp_11 = (temp_10[13:0] - temp_1);
    assign temp_12 = $unsigned(((((((temp_10 - temp_9) ^ temp_6[1:1]) ^ temp_7) * temp_10[14:6]) * input_data) | temp_0[6:5]));
    assign temp_13 = $unsigned(temp_0);
    assign temp_14 = (((((temp_6 - temp_1) - temp_6) * temp_6) - temp_8[13:0]) ^ temp_12);
    assign temp_15 = (temp_5[2:0] - temp_8[18:11]);
    assign temp_16 = temp_5 ? $unsigned(((((((temp_1 ^ input_data) - temp_1) * temp_15[7:0]) | temp_10) + temp_11) | temp_12)) : $signed(temp_10);
    assign temp_17 = $signed((temp_0[6:1] ^ temp_13));
    assign temp_18 = temp_7 ? $signed(($signed((($unsigned(((temp_4[5:5] * temp_10) | temp_11)) * temp_6) - temp_4[5:3])) + temp_4)) : $unsigned((((((temp_13[6:0] ^ (~temp_13)) & temp_6) - temp_0) ^ temp_6) << temp_3));

    assign output_data = ($unsigned((((temp_8 * temp_18) - temp_14) | temp_17)) ^ temp_14);

endmodule