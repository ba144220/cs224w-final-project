module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;
    logic [1:0] temp_17;

    assign temp_0 = ($unsigned((input_data + input_data)) - input_data);
    assign temp_1 = ((((input_data | temp_0) + temp_0) ^ temp_0) & temp_0);
    assign temp_2 = ($signed(temp_0[6:0]) + input_data);
    assign temp_3 = $signed((($signed(((temp_1 * temp_0) | temp_1)) + temp_2) + temp_2));
    assign temp_4 = $unsigned((((input_data + temp_1) * temp_2) ^ input_data));
    assign temp_5 = ((input_data | temp_2) * input_data);
    assign temp_6 = ($unsigned(temp_3) + temp_1[9:0]);
    assign temp_7 = {19'b0, ($unsigned(temp_4) | temp_0[5:0])};
    assign temp_8 = ((((temp_1[18:0] & temp_4) + temp_5) + temp_3) | temp_2);
    assign temp_9 = temp_7;
    assign temp_10 = (temp_9 & temp_9);
    assign temp_11 = ($unsigned((temp_9[3:0] - temp_5)) + temp_2);
    assign temp_12 = ((temp_9 + temp_1) ^ temp_11);
    assign temp_13 = ($signed((($unsigned((temp_6 & temp_0)) * temp_6) * temp_4)) & temp_12[8:0]);
    assign temp_14 = ((((temp_1 + temp_0) - temp_10) * temp_11) * temp_1);
    assign temp_15 = (temp_14 - temp_1);
    assign temp_16 = (((temp_12 | temp_3) & temp_1) | temp_15);
    assign temp_17 = $unsigned(temp_11);

    assign output_data = temp_4;

endmodule