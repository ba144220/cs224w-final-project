module top (
    input [3:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;

    assign temp_0 = ((((((input_data | input_data) + input_data) + (~input_data)) ^ input_data) + input_data) | input_data);
    assign temp_1 = (temp_0 - temp_0[24:17]);
    assign temp_2 = (((temp_1 - input_data) * temp_1) & (~temp_1));
    assign temp_3 = ((($unsigned(($unsigned((temp_0[24:1] - temp_2)) + temp_1)) | temp_1) & input_data[2:0]) - input_data[2:0]);
    assign temp_4 = (((temp_0 + temp_3) ^ temp_1) * temp_0);
    assign temp_5 = (((((temp_2 * temp_0) * temp_3) ^ temp_4) | input_data) & input_data);
    assign temp_6 = ((((((((((input_data - (~temp_4)) + (~temp_5)) - temp_1[8:8]) * input_data) * input_data) * input_data) * (~temp_5)) ^ temp_3) + temp_1) + temp_5);
    assign temp_7 = temp_0 ? ((temp_1[8:8] | temp_2) * temp_5) : ($signed((((($unsigned(((temp_5 | temp_1) & temp_3)) & temp_4) - (~temp_6)) | (~temp_4)) * temp_3)) * temp_3);
    assign temp_8 = temp_5 ? ((temp_7 * temp_4) & input_data) : ($signed(((((((temp_2 + temp_4) - input_data) * temp_0) + temp_3) + input_data) ^ input_data)) - temp_5);
    assign temp_9 = (((((temp_4 | (~temp_3)) ^ input_data[2:1]) - temp_1) & input_data[2:1]) & temp_8);
    assign temp_10 = (((temp_1 - temp_9[1:1]) + temp_7[13:6]) - temp_0);
    assign temp_11 = (temp_0 + temp_5);
    assign temp_12 = temp_8;
    assign temp_13 = (((((((temp_1 ^ temp_5) & temp_4) | temp_6) ^ input_data) | (~temp_1)) + temp_11) & (~temp_5));
    assign temp_14 = (temp_7 + temp_6);
    assign temp_15 = ((((((((((temp_11 * temp_13) + temp_5) | temp_6) | temp_2) * (~temp_8)) & temp_6) | temp_0) ^ (~temp_11)) & temp_0[24:4]) * (~temp_5));

    assign output_data = $signed((((((((($signed(temp_13[24:14]) * temp_4) & temp_5) ^ (~temp_9)) + temp_9) - temp_1) ^ temp_8) - temp_11) ^ temp_10));

endmodule