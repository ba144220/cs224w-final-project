module top (
    input [5:0] input_data,
    output [9:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;

    assign temp_0 = $signed(input_data);
    assign temp_1 = ($unsigned(temp_0[4:0]) * temp_0[3:0]);
    assign temp_2 = (temp_0[4:0] ^ input_data);
    assign temp_3 = $unsigned(($signed((temp_2 - input_data)) | temp_0[2:0]));
    assign temp_4 = ($signed(input_data) >= temp_0);
    logic [6:0] expr_554950;
    assign expr_554950 = ($signed(temp_1[2:0]) + temp_4);
    assign temp_5 = temp_1 ? expr_554950[4:0] : $signed(($signed(input_data[4:0]) & temp_0));
    assign temp_6 = temp_2;
    logic [31:0] expr_942638;
    assign expr_942638 = ($unsigned(($signed(temp_1) - temp_5)) ^ temp_2);
    assign temp_7 = expr_942638[25:0];
    assign temp_8 = ($signed(temp_7) << temp_0);
    assign temp_9 = temp_5;
    assign temp_10 = temp_4;
    assign temp_11 = temp_8;
    assign temp_12 = ($signed(temp_5) >> temp_3);
    assign temp_13 = $signed(($unsigned(temp_0[6:3]) + temp_7));
    assign temp_14 = temp_7;
    assign temp_15 = ($unsigned(($unsigned(temp_5) << temp_2)) ^ temp_14[4:0]);

    assign output_data = (($unsigned(temp_2) + temp_5) + temp_5);

endmodule