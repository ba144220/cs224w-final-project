module top (
    input [9:0] input_data,
    output [39:0] output_data
);

    logic [23:0] temp_0;
    logic [17:0] temp_1;
    logic [8:0] temp_2;
    logic [11:0] temp_3;
    logic [0:0] temp_4;
    logic [21:0] temp_5;
    logic [29:0] temp_6;
    logic [5:0] temp_7;
    logic [21:0] temp_8;
    logic [2:0] temp_9;
    logic [24:0] temp_10;
    logic [10:0] temp_11;
    logic [28:0] temp_12;
    logic [27:0] temp_13;
    logic [10:0] temp_14;
    logic [10:0] temp_15;
    logic [15:0] temp_16;
    logic [3:0] temp_17;

    assign temp_0 = input_data[9:9] ? input_data : ($unsigned(24'd7042744) & input_data);
    assign temp_1 = input_data;
    assign temp_2 = ($unsigned(temp_0) | input_data[9:1]);
    logic [23:0] expr_910856;
    assign expr_910856 = temp_0;
    assign temp_3 = expr_910856[11:0];
    assign temp_4 = (input_data[8:8] | temp_0);
    assign temp_5 = ($signed(($unsigned((($signed(($signed(temp_3) | temp_0)) <= input_data) - input_data)) * temp_1)) | input_data);
    assign temp_6 = ($signed((temp_0 + temp_3)) - (~temp_2));
    assign temp_7 = input_data[8:3];
    assign temp_8 = (($signed(($unsigned(temp_4) + (~temp_6))) ^ temp_4) + temp_0[23:8]);
    assign temp_9 = $unsigned(($signed(temp_6) - temp_2[1:0]));
    assign temp_10 = temp_6;
    assign temp_11 = ($unsigned(temp_1[3:0]) * temp_0);
    assign temp_12 = ($signed((($signed(input_data) + (~input_data)) * temp_0)) + input_data);
    assign temp_13 = ($signed((($unsigned(temp_7) >> temp_5) ^ temp_2)) << temp_8);
    assign temp_14 = ((($signed(($unsigned(temp_8) * temp_2)) & temp_9) * temp_9) + temp_0);
    assign temp_15 = (((($unsigned(temp_5) ^ temp_8) + temp_5) - temp_9) ^ temp_5[13:0]);
    assign temp_16 = temp_2 ? ($signed(temp_0) ^ temp_5[19:0]) : (($unsigned(temp_7) + temp_4) << (~temp_4));
    assign temp_17 = ($signed((($signed(($unsigned(($unsigned(temp_16) * (~temp_6))) + temp_3)) * temp_11) - temp_6[27:0])) * temp_2);

    assign output_data = ($signed((($unsigned((($signed(temp_11) & temp_1) | temp_13)) ^ temp_7) | temp_5[4:0])) & temp_15[7:0]);

endmodule