module top (
    input [11:0] input_data,
    output [16:0] output_data
);

    logic [22:0] temp_0;
    logic [1:0] temp_1;
    logic [29:0] temp_2;
    logic [15:0] temp_3;
    logic [3:0] temp_4;
    logic [10:0] temp_5;
    logic [7:0] temp_6;
    logic [23:0] temp_7;
    logic [30:0] temp_8;
    logic [15:0] temp_9;
    logic [24:0] temp_10;
    logic [6:0] temp_11;
    logic [15:0] temp_12;
    logic [0:0] temp_13;
    logic [13:0] temp_14;
    logic [26:0] temp_15;
    logic [17:0] temp_16;

    assign temp_0 = input_data[6:6] ? (input_data * input_data) : ((input_data - input_data) * 23'd2444472);
    logic [27:0] expr_289067;
    assign expr_289067 = (((((input_data[6:5] - temp_0) & (~temp_0)) - input_data[2:1]) & temp_0) * 2'd0);
    assign temp_1 = expr_289067[1:0];
    assign temp_2 = ((((temp_0 | input_data) < (~temp_1)) == temp_1) * input_data);
    assign temp_3 = input_data[2:2] ? ((((input_data & temp_0) & input_data) | temp_1) ^ input_data) : (((((temp_1 * input_data) ^ input_data) * input_data) & temp_0) | temp_1);
    assign temp_4 = ((((input_data[3:0] & input_data[5:2]) & (~temp_0)) - temp_2) + input_data[3:0]);
    logic [17:0] expr_660032;
    assign expr_660032 = ((temp_4 - temp_3) * input_data[11:1]);
    assign temp_5 = expr_660032[10:0];
    assign temp_6 = ((((temp_2 & input_data[11:4]) * temp_3) - (~temp_0)) - 8'd140);
    assign temp_7 = (((((temp_3 ^ -24'd2368503) * 24'd4445278) & temp_0) & temp_5) & temp_5);
    assign temp_8 = (((temp_4 | input_data) + temp_3) * temp_1);
    assign temp_9 = (((((temp_7 & 16'd14183) * temp_1) * (~temp_7)) ^ temp_8) + temp_4);
    assign temp_10 = (temp_0 | temp_6);
    assign temp_11 = temp_6 ? temp_3 : ((temp_6 ^ temp_10) | temp_2);
    assign temp_12 = ((input_data ^ temp_1) > temp_4);
    assign temp_13 = ((temp_7 - temp_5) & temp_9);
    assign temp_14 = ((temp_12 + temp_6) == temp_0);
    assign temp_15 = (((temp_10 + (~temp_13)) & temp_8) - temp_14);
    assign temp_16 = (((temp_9 - temp_4) * temp_2) ^ temp_1);

    assign output_data = temp_10 ? temp_4 : temp_8;

endmodule