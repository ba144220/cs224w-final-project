module top (
    input [2:0] input_data,
    output [2:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;

    assign temp_0 = $signed(((input_data + input_data) & input_data));
    assign temp_1 = ((input_data | temp_0) | temp_0);
    assign temp_2 = ((temp_0 - input_data) ^ input_data);
    assign temp_3 = {14'b0, temp_0};
    assign temp_4 = {4'b0, (($unsigned(temp_2) + (~temp_0[3:0])) - temp_0)};
    assign temp_5 = $signed(temp_4);
    assign temp_6 = $unsigned(((temp_4 - temp_5) - temp_3));
    assign temp_7 = $unsigned(temp_1[21:0]);
    assign temp_8 = temp_7[2:0] ? ($unsigned(($unsigned(temp_5) | (~temp_2[7:0]))) + temp_2) : ((temp_6[2:1] & (~temp_2)) + temp_4);
    assign temp_9 = $signed(((temp_7 | (~temp_4[10:0])) & temp_5));

    assign output_data = ((temp_1[22:0] & temp_0) * temp_4);

endmodule