module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;

    assign temp_0 = ($unsigned((input_data + input_data)) * input_data);
    assign temp_1 = input_data;
    assign temp_2 = (temp_0 + temp_1);
    assign temp_3 = ($signed(($signed((temp_0 * temp_0[6:1])) | temp_0)) + input_data);
    assign temp_4 = $unsigned(temp_1);
    assign temp_5 = ($unsigned((temp_0 - temp_0)) + temp_4);
    assign temp_6 = ($signed(temp_3) - temp_0[3:0]);
    assign temp_7 = input_data[4:4] ? ($unsigned((($signed(temp_5) + temp_6) ^ temp_3)) & (~26'd25670156)) : $signed(temp_3);
    assign temp_8 = temp_1 ? ((($unsigned(temp_3) | (~temp_7)) | temp_2[3:0]) + temp_5[4:4]) : ($signed(((temp_5 ^ temp_1) & temp_2)) * temp_0[6:3]);
    assign temp_9 = (((temp_0 * temp_7) & temp_7) * temp_1);

    assign output_data = $unsigned(temp_2);

endmodule