module top (
    input [6:0] input_data,
    output [5:0] output_data
);

    logic [31:0] temp_0;
    logic [16:0] temp_1;
    logic [2:0] temp_2;
    logic [0:0] temp_3;
    logic [9:0] temp_4;
    logic [30:0] temp_5;
    logic [23:0] temp_6;
    logic [20:0] temp_7;
    logic [1:0] temp_8;
    logic [17:0] temp_9;
    logic [31:0] temp_10;
    logic [12:0] temp_11;
    logic [26:0] temp_12;
    logic [6:0] temp_13;

    assign temp_0 = ($signed(($unsigned(input_data) * input_data)) + input_data);
    assign temp_1 = $unsigned(($signed(temp_0) & temp_0[29:0]));
    assign temp_2 = ($unsigned(temp_0[31:11]) | input_data[4:2]);
    assign temp_3 = ($signed(($signed(($unsigned(input_data[4:4]) ^ input_data[6:6])) & temp_1)) - temp_2);
    assign temp_4 = ($unsigned(($unsigned((temp_3 & temp_3)) & temp_2)) * temp_3);
    assign temp_5 = temp_0;
    assign temp_6 = temp_1;
    assign temp_7 = ($unsigned(($signed(($signed(temp_5) + temp_5)) ^ temp_1)) ^ (~temp_6));
    assign temp_8 = ($signed(($signed(($signed(temp_3) | (~temp_2[2:1]))) ^ (~temp_6))) | input_data[6:5]);
    assign temp_9 = ($signed(temp_2) | temp_6);
    assign temp_10 = ($signed(temp_2) ^ temp_1[2:0]);
    assign temp_11 = $signed(temp_9);
    assign temp_12 = ($unsigned(($unsigned(($unsigned(27'd114173553) ^ temp_4)) - temp_0)) ^ temp_8[1:0]);
    assign temp_13 = ($unsigned(($signed(temp_2[2:0]) + temp_7)) & temp_3);

    logic [26:0] expr_168261;
    assign expr_168261 = temp_12;
    assign output_data = expr_168261[5:0];

endmodule