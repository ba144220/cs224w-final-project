module top (
    input [2:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;
    logic [25:0] temp_16;

    assign temp_0 = ($signed(($unsigned(($unsigned(input_data) & input_data)) & input_data)) ^ input_data);
    assign temp_1 = ($signed((($unsigned(($signed(($unsigned(($signed(($unsigned(($unsigned(($signed((($signed((($unsigned(input_data) & temp_0) | temp_0)) | input_data) * temp_0)) & temp_0)) * input_data)) + temp_0[24:22])) | temp_0)) | temp_0)) | temp_0)) & input_data) - input_data)) & input_data);
    assign temp_2 = temp_0;
    assign temp_3 = (($unsigned((($unsigned(input_data) - temp_0) | temp_1)) * temp_2) ^ temp_2);
    assign temp_4 = ($unsigned(($signed((($unsigned(($unsigned(((((($unsigned((($signed(($unsigned(temp_2) | input_data)) ^ temp_2) | temp_1)) ^ temp_3) + temp_3) | temp_0[24:3]) * input_data) * temp_2)) | temp_1)) | temp_2) ^ temp_1)) & temp_0)) - temp_3);
    assign temp_5 = (($signed(($signed(($signed(($unsigned(temp_2) - temp_3)) | temp_1)) * (~temp_0))) - 9'd459) & (~temp_4));
    assign temp_6 = (($signed(($signed(($unsigned((temp_1 | temp_2)) ^ temp_5)) & temp_4)) * temp_2) + temp_5);
    assign temp_7 = (($signed(($unsigned((($signed(($unsigned(($signed(($signed(($signed(temp_1) + temp_6)) - (~14'd6941))) + temp_4)) + temp_6)) ^ input_data) ^ input_data)) + temp_5)) - (~temp_3)) - temp_5);
    assign temp_8 = (($unsigned((($signed(($signed(($signed((($signed(($signed(($signed((input_data & input_data)) - temp_5)) | input_data)) | temp_3) * temp_6)) + temp_3[2:2])) | temp_0)) + temp_5) * temp_0)) | input_data) & temp_2);
    assign temp_9 = ($signed((($signed(($signed(($unsigned(($signed((($unsigned(temp_2) * temp_0) ^ input_data[2:1])) | temp_1)) - (~temp_5))) * temp_8)) * input_data[2:1]) - temp_2)) & temp_6);
    assign temp_10 = (($unsigned(((($unsigned(($signed((($unsigned(input_data) * input_data) ^ temp_3[2:1])) - temp_7)) + (~temp_7)) | temp_0) ^ temp_5)) + temp_0) * temp_8);
    assign temp_11 = ($unsigned((($signed(($signed((($signed(($signed(($unsigned(($signed(($unsigned(temp_6) - input_data)) | temp_10)) | temp_9)) + temp_0)) ^ temp_4) - temp_10)) | (~temp_0))) & (~temp_10)) ^ temp_5)) | temp_3);
    logic [35:0] expr_645483;
    assign expr_645483 = $unsigned(((($signed(($signed((($signed((($unsigned(($unsigned(($unsigned(($unsigned((temp_7 + input_data)) & temp_3)) & temp_7)) - temp_2)) | temp_1) + temp_8)) ^ temp_10) ^ temp_9)) + temp_7)) & temp_8) ^ temp_0) & temp_0));
    assign temp_12 = expr_645483[29:0];
    assign temp_13 = ((temp_10[29:9] * temp_5) - temp_1);
    assign temp_14 = ($signed(($signed(($unsigned((($unsigned(($unsigned((($signed(($unsigned(($signed(temp_6) & temp_10)) * temp_0)) - temp_0) * temp_5)) * (~temp_2))) - temp_8) * temp_13)) | temp_6)) - temp_7)) - temp_6);
    assign temp_15 = ($unsigned(($unsigned(($signed(($signed((($unsigned(((($unsigned(($signed(temp_14) * temp_5)) + temp_4) - temp_13) | input_data)) - temp_1) & temp_7)) & temp_6)) * temp_1)) | temp_3)) - (~temp_8));
    assign temp_16 = $unsigned((($unsigned(temp_11) + temp_10) - temp_12));

    assign output_data = {8'b0, ($signed(temp_3) ^ temp_3)};

endmodule