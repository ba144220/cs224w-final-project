module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;

    assign temp_0 = (((((($signed((input_data & input_data)) - input_data) | input_data) & input_data) & input_data) | input_data) * input_data);
    assign temp_1 = $signed((($signed(($signed(($signed(($signed(((input_data & temp_0) | input_data)) - input_data)) + input_data)) & input_data)) + temp_0[1:0]) ^ temp_0));
    assign temp_2 = $unsigned(($unsigned(temp_0) | input_data));
    assign temp_3 = (($signed(($unsigned(($signed(((input_data | input_data) - temp_0)) + input_data)) | input_data)) & temp_0) + temp_2);
    logic [23:0] expr_691179;
    assign expr_691179 = ((($unsigned((((temp_3 - temp_3) | temp_2) & (~input_data))) >> (~temp_0[1:0])) >> temp_2) - temp_0[3:0]);
    assign temp_4 = expr_691179[16:0];
    assign temp_5 = temp_3[12:0];
    assign temp_6 = (($unsigned((($signed(((temp_1[20:0] * temp_5) + (~temp_1))) + input_data) ^ input_data)) | input_data) * temp_1);
    assign temp_7 = (((($signed((((temp_5 & temp_2) | temp_5) | temp_3)) * temp_5) - temp_4) | temp_1) | temp_4);
    assign temp_8 = ($unsigned((($signed((($signed(temp_1) == input_data) * temp_6)) + temp_6) + temp_6)) * temp_4[11:0]);
    assign temp_9 = ($signed(temp_2) * temp_7);
    assign temp_10 = ($signed(((($signed(($signed(temp_7) - temp_7)) & temp_5) & temp_5) ^ temp_6)) ^ temp_9);

    assign output_data = ($signed((temp_0[2:0] * temp_1)) | temp_5);

endmodule