module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;

    assign temp_0 = input_data;
    assign temp_1 = ($unsigned((temp_0 * input_data)) ^ input_data);
    assign temp_2 = ($signed(($signed((($unsigned(($unsigned((($unsigned(temp_1) | temp_1) | temp_1)) | temp_1)) + temp_1) ^ temp_0)) * temp_0[5:1])) + temp_0[1:0]);
    assign temp_3 = temp_0[5:3] ? (($signed((($signed(($unsigned(((((temp_1[15:0] | temp_2[5:0]) ^ temp_0) - temp_1) * temp_1)) * temp_0)) + input_data) | temp_1)) & temp_0[5:1]) - temp_2) : ($signed(((($signed(($signed(($signed(($signed((($signed(($signed(($unsigned(temp_2) | temp_0)) * temp_1)) ^ input_data) | temp_0)) & temp_2)) * temp_0)) | temp_0)) * temp_1) & temp_1) + temp_2)) & input_data);
    assign temp_4 = ((($unsigned(((($unsigned(($signed((input_data + temp_1)) ^ temp_2)) | temp_1[23:9]) ^ temp_2) ^ temp_1)) + temp_3) | temp_1[23:18]) ^ input_data);
    assign temp_5 = ($signed(($signed(($signed(($signed(($unsigned(($signed((($signed((input_data + input_data)) == input_data) * temp_3)) + temp_3)) + temp_4)) * temp_4)) | temp_3)) * temp_0)) - temp_3);
    assign temp_6 = ($unsigned(($signed(temp_2[10:4]) & temp_5)) | temp_3);
    assign temp_7 = $signed((($signed(($signed(($signed((($signed(input_data) | temp_5) & temp_1)) - temp_5)) & temp_3[19:11])) - temp_1) | temp_2));
    assign temp_8 = ($unsigned((($signed((($signed(($signed(($signed(($signed(($unsigned(temp_6[2:2]) & temp_5)) & input_data)) + temp_2)) & temp_0)) + temp_7[8:0]) - temp_0[5:0])) | temp_3) - temp_3)) ^ temp_2);
    assign temp_9 = ($signed((temp_8 | temp_4)) + temp_3);
    assign temp_10 = ($signed(($unsigned(($signed(($signed((($signed((($unsigned(($signed((($unsigned(temp_9) + temp_8) ^ temp_3)) | temp_6)) ^ temp_4[16:14]) | temp_3[19:6])) & temp_6) & temp_5[13:10])) | temp_9)) * temp_0)) * temp_1)) - temp_6);
    assign temp_11 = (($unsigned(($signed((($signed(($unsigned(($unsigned(($signed(($signed(temp_3) * temp_6)) - temp_6[2:2])) - temp_0)) + temp_6)) & temp_7) - temp_3)) + temp_8)) ^ temp_0) + temp_5);

    assign output_data = temp_10[22:0];

endmodule