module top (
    input [3:0] input_data,
    output [37:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;
    logic [14:0] temp_13;
    logic [9:0] temp_14;

    assign temp_0 = ((((input_data + input_data) << input_data) >> input_data) * input_data);
    assign temp_1 = {12'b0, $unsigned((((temp_0 + input_data) | input_data) * temp_0))};
    assign temp_2 = (((temp_0 | temp_0[8:1]) | temp_0) * input_data);
    assign temp_3 = ($signed((((temp_1 * temp_0) | temp_0) | (~temp_2))) * temp_1);
    assign temp_4 = temp_1;
    assign temp_5 = (((temp_2 * temp_1) & temp_4) ^ temp_3);
    assign temp_6 = $unsigned(($unsigned(($signed((input_data & temp_3)) ^ (~input_data))) & input_data));
    assign temp_7 = (((($unsigned(input_data) * temp_0) - temp_0) - temp_4) + (~temp_0[8:1]));
    assign temp_8 = $unsigned(($unsigned(($signed(temp_4) + temp_0)) | temp_6[16:14]));
    assign temp_9 = temp_4 ? (((temp_5 * temp_1) & temp_5[30:19]) - temp_0) : $unsigned(temp_4);
    assign temp_10 = temp_8;
    assign temp_11 = (temp_4 * temp_1);
    assign temp_12 = $signed(((((temp_10 - temp_11) - temp_3) | temp_4) * temp_4));
    assign temp_13 = ((($unsigned(temp_10) ^ temp_6) ^ temp_10) * temp_9);
    assign temp_14 = {1'b0, temp_0};

    assign output_data = $unsigned(((($signed(temp_10) << temp_2[30:9]) | temp_1) >> temp_4));

endmodule