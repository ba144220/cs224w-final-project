module top (
    input [7:0] input_data,
    output [9:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;
    logic [26:0] temp_10;
    logic [4:0] temp_11;

    assign temp_0 = $signed(($signed(((((($unsigned(((input_data ^ input_data) - 26'd38870700)) | (~input_data)) + input_data) & input_data) & input_data) - input_data)) ^ input_data));
    assign temp_1 = $unsigned(((($signed(($signed(($signed(($unsigned(((temp_0 & (~temp_0)) ^ (~temp_0))) & temp_0)) & temp_0)) ^ (~temp_0))) ^ temp_0) | temp_0) + temp_0));
    assign temp_2 = temp_0[5:0] ? $signed((((((($unsigned((($unsigned(temp_0) * input_data[7:3]) & temp_1[1:0])) & input_data[4:0]) ^ (~temp_0)) * temp_0) ^ temp_0) | temp_0) | input_data[6:2])) : ($unsigned(((temp_0 ^ temp_0) - temp_1[3:0])) + input_data[5:1]);
    assign temp_3 = ((($signed(((((temp_0[24:0] ^ temp_2) - temp_0) & 7'd117) | (~temp_2[2:0]))) & input_data[6:0]) | (~temp_2)) | temp_0);
    assign temp_4 = ($unsigned(($unsigned((($unsigned((($unsigned(((temp_3 | input_data) - input_data)) ^ temp_0) ^ temp_1)) + temp_3) & temp_1)) & (~temp_0))) - (~input_data));
    assign temp_5 = $unsigned(((((temp_3 + temp_1) * temp_1[1:0]) | temp_2) - temp_1));
    assign temp_6 = temp_4;
    assign temp_7 = temp_3 ? $unsigned(($unsigned(($signed((($signed(($unsigned(($signed(temp_1) ^ (~temp_1))) ^ input_data[2:0])) ^ (~input_data[7:5])) & temp_2)) * temp_1[2:0])) - temp_0[3:0])) : (($signed(((($signed((((input_data[6:4] & temp_5) + temp_5) - input_data[6:4])) ^ (~temp_5)) * input_data[5:3]) ^ temp_1[3:1])) | temp_4[16:0]) ^ temp_1);
    assign temp_8 = ((($signed(temp_4) > temp_4) | temp_7) - 6'd57);
    assign temp_9 = temp_8 ? $unsigned(((((($signed((((temp_7 + temp_7) & (~temp_5[2:0])) - temp_4)) + temp_6) ^ temp_3) & temp_6) + temp_6) + temp_8[4:0])) : ($signed((($unsigned(((($unsigned(temp_6[11:0]) - temp_8) & (~temp_8)) - temp_3)) | (~temp_4)) | temp_3[2:0])) & input_data);
    assign temp_10 = (temp_7 + temp_2);
    assign temp_11 = ($unsigned((((((((temp_9 | (~temp_10)) - (~temp_9)) | temp_4) & (~temp_0)) >> temp_10) & (~temp_5)) | temp_8[4:0])) & temp_3);

    assign output_data = temp_6[1:0];

endmodule