module top (
    input [5:0] input_data,
    output [9:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;

    assign temp_0 = ($signed(($signed(($unsigned((input_data - input_data)) * input_data)) * 7'd99)) + input_data);
    assign temp_1 = ($signed(($signed((temp_0 + (~temp_0))) ^ temp_0)) | temp_0);
    assign temp_2 = {4'b0, ($unsigned(temp_0) ^ temp_1)};
    assign temp_3 = $signed(($unsigned((($signed(temp_0[6:1]) & temp_1) + temp_0)) | temp_0[6:5]));
    assign temp_4 = $signed((input_data - temp_2));
    assign temp_5 = input_data[4:0];
    assign temp_6 = temp_4 ? $unsigned(($unsigned(($signed(input_data[4:3]) | temp_5)) * input_data[1:0])) : ($unsigned((($unsigned(((temp_3[9:3] + temp_2) | temp_1)) & input_data[1:0]) * temp_1[25:17])) * temp_0);
    assign temp_7 = temp_4;
    assign temp_8 = $unsigned(($unsigned(temp_1) - (~temp_2)));
    assign temp_9 = $signed(($unsigned(($unsigned(($unsigned(($signed(($unsigned(temp_6) - temp_0)) | temp_8)) * temp_5[4:2])) * temp_5)) * temp_5));

    logic [31:0] expr_536143;
    assign expr_536143 = ($unsigned(($signed(($signed((temp_1 & temp_9)) & temp_7)) >> temp_6)) | temp_2);
    assign output_data = temp_2 ? expr_536143[9:0] : $signed(temp_5);

endmodule