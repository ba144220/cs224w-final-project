module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;
    logic [1:0] temp_17;

    assign temp_0 = ($unsigned((($unsigned((($signed(($unsigned(input_data) ^ input_data)) | input_data) | input_data)) * input_data) - (~input_data))) + input_data);
    assign temp_1 = ($unsigned(temp_0) | temp_0[6:2]);
    assign temp_2 = $signed(input_data);
    assign temp_3 = ($unsigned(($signed(($signed(10'd909) * temp_1)) * input_data)) - temp_0[2:0]);
    assign temp_4 = input_data;
    assign temp_5 = ((($unsigned(temp_3) + (~temp_2)) + input_data[4:0]) ^ temp_0[6:2]);
    logic [8:0] expr_967166;
    assign expr_967166 = ($unsigned(((input_data[3:2] * input_data[1:0]) ^ temp_0)) + input_data[4:3]);
    assign temp_6 = expr_967166[1:0];
    assign temp_7 = ($signed((($unsigned((input_data | temp_1)) & input_data) * temp_1[3:0])) + temp_2[30:18]);
    assign temp_8 = ($signed(($signed(($unsigned(temp_5) != temp_1)) - input_data)) ^ temp_0[6:3]);
    assign temp_9 = ($unsigned(($unsigned((temp_0 * temp_7)) & temp_7)) & temp_2);
    assign temp_10 = $signed(temp_5);
    assign temp_11 = (($unsigned(($signed(($unsigned(($unsigned(($signed(temp_2) | 24'd3919974)) - temp_10)) ^ temp_5)) & temp_5)) ^ temp_5) ^ input_data);
    assign temp_12 = ($signed(($unsigned(($unsigned(($signed(temp_4[5:4]) | temp_8)) - temp_5[3:0])) ^ (~temp_11))) * temp_11);
    assign temp_13 = ($unsigned(($unsigned(temp_6) & (~input_data))) + temp_0);
    assign temp_14 = $unsigned(($signed(((($signed((temp_13 & temp_5)) + temp_3) ^ temp_12) ^ 7'd121)) + temp_0));
    assign temp_15 = temp_13[4:0];
    assign temp_16 = ($signed(($signed((($unsigned(($signed(temp_6) ^ temp_9)) - temp_9) & temp_13)) << temp_6)) * temp_10[13:0]);
    assign temp_17 = $signed((($signed(($unsigned(temp_6) + (~temp_10))) - temp_0) ^ (~temp_11)));

    assign output_data = (($unsigned(($signed(($signed(($signed(temp_15) - temp_12)) + temp_1)) | temp_11)) - temp_17[1:1]) | temp_15);

endmodule