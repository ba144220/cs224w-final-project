module top (
    input [5:0] input_data,
    output [37:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;
    logic [14:0] temp_13;
    logic [9:0] temp_14;
    logic [24:0] temp_15;
    logic [0:0] temp_16;
    logic [4:0] temp_17;

    logic [11:0] expr_113371;
    assign expr_113371 = $signed(($unsigned(($signed(($unsigned(($unsigned(($signed(($unsigned(($unsigned(($signed(($unsigned(input_data) > input_data)) >= input_data)) & input_data)) < input_data)) + input_data)) >= input_data)) - 9'd495)) * 9'd425)) + input_data));
    assign temp_0 = expr_113371[8:0];
    assign temp_1 = $unsigned(temp_0[8:6]);
    assign temp_2 = $unsigned(($unsigned((($signed((($unsigned(($signed(($unsigned(input_data) | input_data)) * temp_1)) + temp_0[6:0]) ^ (~temp_1[2:0]))) * temp_1) | temp_1[1:0])) - temp_0));
    assign temp_3 = $unsigned(($unsigned(($signed(($unsigned(temp_1) | temp_0[8:4])) * temp_2[20:0])) * temp_2));
    assign temp_4 = ($signed(($signed(($unsigned(($unsigned(($signed((1'd1 | (~temp_1))) - temp_1)) - temp_1)) * temp_3[4:2])) - temp_2)) & temp_2);
    assign temp_5 = input_data;
    assign temp_6 = ($unsigned(temp_2) & (~temp_4));
    assign temp_7 = ($signed(($unsigned(($unsigned(($unsigned((($unsigned(($signed(($unsigned(($unsigned(($unsigned(temp_2) * (~temp_5[30:7]))) & temp_1)) * temp_5)) ^ temp_2)) & temp_0) + temp_0)) + (~temp_6))) | temp_2)) & temp_6)) + temp_1);
    assign temp_8 = $unsigned(($signed(($signed(($signed(($signed(($signed(($unsigned(($unsigned(input_data) ^ temp_7)) | temp_3)) | input_data)) & temp_5)) ^ temp_7)) + input_data)) ^ temp_1));
    assign temp_9 = $unsigned(($unsigned(($unsigned(($unsigned(($signed(temp_1) - (~temp_4))) ^ temp_7[11:0])) ^ temp_4)) ^ temp_5));
    assign temp_10 = ($signed((($unsigned(($signed(($unsigned(($unsigned(($unsigned(($signed(temp_0) | temp_2)) - input_data)) * temp_1[6:0])) * temp_4)) | temp_5)) + (~temp_9[4:0])) ^ (~temp_6))) | temp_6);
    assign temp_11 = $signed(($signed(($unsigned(($signed(($unsigned(($signed(($unsigned(($unsigned(temp_8) & (~input_data))) - temp_0[4:0])) - temp_3[4:0])) - temp_1[23:12])) + input_data)) | temp_0)) - temp_3));
    assign temp_12 = ($signed(($unsigned(($signed(($signed(($signed(($unsigned(temp_7) - temp_0)) - input_data)) - (~temp_0))) - (~temp_2[1:0]))) ^ temp_6[16:0])) + (~temp_3));
    logic [19:0] expr_180015;
    assign expr_180015 = ($unsigned(($signed(($signed(($unsigned(($signed(($signed(($unsigned(temp_8) ^ input_data)) + temp_10[6:0])) | temp_3)) ^ temp_4)) & temp_6)) ^ temp_8)) ^ temp_4);
    assign temp_13 = expr_180015[14:0];
    assign temp_14 = temp_10[8:0];
    assign temp_15 = ($signed(($signed(($unsigned(($unsigned(($signed(($signed(($signed((($signed(temp_11) + temp_6) ^ temp_11[5:0])) + temp_4)) | temp_14)) + temp_13)) - temp_10)) | temp_12)) | (~temp_4))) | temp_5);
    assign temp_16 = ($signed(temp_6) ^ temp_13);
    assign temp_17 = $unsigned(temp_3[2:0]);

    assign output_data = $signed(($unsigned(($signed(($signed(temp_11) * temp_4)) ^ temp_9)) * temp_14));

endmodule