module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;

    assign temp_0 = $unsigned(input_data);
    assign temp_1 = ($unsigned(($signed(($unsigned(temp_0) - input_data)) | temp_0)) & temp_0);
    assign temp_2 = ($signed(($signed(($signed(($signed(($signed((($unsigned(temp_0) & temp_1) + input_data)) ^ temp_0)) * temp_0[5:1])) + temp_0[1:0])) ^ temp_0[5:2])) | input_data);
    assign temp_3 = $unsigned(($signed(($unsigned(($signed(($unsigned(($unsigned(($signed(temp_0[3:0]) + temp_0)) * temp_2)) * temp_0)) + input_data)) | input_data)) & temp_0[5:1]));
    assign temp_4 = $signed(($unsigned(($unsigned(($unsigned(($unsigned((($unsigned(input_data) & temp_0) & temp_0)) + input_data)) + 17'd121461)) * temp_2[10:8])) & temp_2[10:2]));
    assign temp_5 = ($signed(($signed(($signed((($unsigned(($unsigned(($signed(temp_2[10:6]) * temp_3)) & temp_3)) ^ 14'd4800) ^ input_data)) ^ input_data)) & temp_4)) - (~temp_2));
    assign temp_6 = ($signed(($unsigned((($signed(($signed(($unsigned((($unsigned(temp_5) & temp_4) - temp_1)) + (~temp_4))) - input_data)) - temp_4) & temp_4)) * temp_3)) * temp_4);
    assign temp_7 = ($unsigned(($signed(input_data) + temp_3)) ^ temp_5[12:0]);
    assign temp_8 = $signed(($unsigned(($signed(($signed(($signed(28'd209984069) | temp_2)) - temp_0[5:4])) * temp_2)) ^ temp_4[16:8]));
    assign temp_9 = ($unsigned(($signed(($signed(($unsigned(($unsigned((($unsigned(($unsigned(temp_5) | temp_5)) ^ temp_1) & temp_2)) - temp_6[2:0])) * temp_2)) * temp_6[2:1])) * input_data)) & temp_2);
    assign temp_10 = ($unsigned(($unsigned(($signed(($signed(($signed((($signed(temp_9) | temp_7) + temp_7[10:9])) * temp_0)) + temp_7[8:0])) - temp_8[7:0])) * temp_3[16:0])) & temp_0);
    assign temp_11 = ($unsigned(($unsigned(temp_3) * temp_6[2:0])) & temp_8);

    assign output_data = temp_8 ? ($unsigned(($unsigned(($unsigned(($signed(($unsigned(($signed(temp_10[9:0]) ^ temp_11[28:25])) * temp_0)) + temp_10)) ^ temp_4)) + temp_7)) + temp_3) : ($unsigned(($signed(temp_7) & temp_7)) | temp_5);

endmodule