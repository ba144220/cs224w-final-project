module top (
    input [3:0] input_data,
    output [31:0] output_data
);

    logic [16:0] temp_0;
    logic [2:0] temp_1;
    logic [0:0] temp_2;
    logic [9:0] temp_3;
    logic [30:0] temp_4;
    logic [23:0] temp_5;
    logic [20:0] temp_6;
    logic [1:0] temp_7;

    assign temp_0 = $unsigned(($unsigned(($signed(($unsigned(input_data) - input_data)) & input_data)) ^ input_data));
    assign temp_1 = (($unsigned((($signed(($unsigned((($unsigned(temp_0) & temp_0[7:0]) - temp_0)) + temp_0[11:0])) * temp_0) & temp_0)) & temp_0) + (~temp_0));
    assign temp_2 = $unsigned(((($unsigned(input_data[3:3]) & temp_1) ^ input_data[1:1]) & input_data[3:3]));
    assign temp_3 = temp_2;
    assign temp_4 = temp_2 ? ($signed(($unsigned(($signed(($unsigned(($signed(($signed(($unsigned(($signed(temp_2) - temp_1[1:0])) ^ input_data)) ^ input_data)) - input_data)) + input_data)) * temp_3)) ^ temp_0)) - temp_2) : ($unsigned(($unsigned(temp_1) | temp_3)) ^ temp_2);
    assign temp_5 = temp_1;
    assign temp_6 = $unsigned(($signed(($signed(temp_0[16:0]) + temp_5)) & temp_4));
    assign temp_7 = (($unsigned(temp_5) ^ temp_3) * temp_2);

    assign output_data = ($unsigned(($unsigned(($unsigned(((($signed(($unsigned(($signed(($unsigned(temp_5) + temp_5)) * temp_0[3:0])) | temp_3)) << temp_7) - temp_2) - temp_2)) >> temp_3)) + temp_5)) & temp_0);

endmodule