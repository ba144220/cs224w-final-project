module top (
    input [3:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;

    assign temp_0 = $signed((($unsigned(((($unsigned(((input_data + input_data) & input_data)) + input_data) + input_data) - input_data)) + input_data) | input_data));
    assign temp_1 = $unsigned((($unsigned(($unsigned(($signed((input_data * temp_0)) ^ input_data)) * temp_0)) - input_data) - input_data));
    assign temp_2 = temp_0 ? ($unsigned(($signed(input_data) - temp_0)) * temp_1) : $signed(((temp_0 & input_data) - input_data));
    assign temp_3 = ((($signed(((($signed((temp_2 ^ input_data[2:0])) < input_data[2:0]) ^ input_data[2:0]) < input_data[3:1])) ^ input_data[2:0]) | temp_1) != temp_2);
    assign temp_4 = (input_data * temp_2);
    assign temp_5 = ($signed(((temp_1 + temp_1) - temp_1)) * 9'd67);
    assign temp_6 = (temp_2 * temp_0);
    assign temp_7 = (temp_1 + temp_6);
    assign temp_8 = $signed((((($signed(((($signed(((temp_2 - temp_7[8:0]) & temp_6)) ^ temp_5) - temp_4) * temp_6)) & temp_5) ^ temp_2) | temp_1) * temp_5[6:0]));

    assign output_data = ($unsigned(($unsigned((($signed((temp_0 ^ temp_5[4:0])) & temp_8) * temp_4)) ^ temp_1)) * temp_7);

endmodule