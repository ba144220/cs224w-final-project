module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;

    assign temp_0 = ((input_data - input_data) * input_data);
    assign temp_1 = $signed(((temp_0 | 26'd41844012) & temp_0));
    assign temp_2 = ((temp_0 ^ temp_1) - input_data);
    assign temp_3 = temp_0;
    assign temp_4 = temp_1 ? $signed(((temp_3 * temp_0) | (~temp_3))) : temp_2;
    assign temp_5 = temp_0;
    assign temp_6 = $signed(temp_1);
    assign temp_7 = $signed(temp_5);
    assign temp_8 = ((temp_7 & temp_4) * input_data);
    assign temp_9 = {2'b0, $unsigned(temp_6)};

    assign output_data = temp_6;

endmodule