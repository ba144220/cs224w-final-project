module top (
    input [3:0] input_data,
    output [36:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;
    logic [0:0] temp_13;
    logic [28:0] temp_14;

    assign temp_0 = (($unsigned((input_data + input_data)) - input_data) | input_data);
    assign temp_1 = ($signed(($signed(($signed(($signed(($signed((($signed(($unsigned(input_data) + input_data)) * input_data) & temp_0)) + (~temp_0))) + temp_0)) | temp_0)) ^ temp_0)) | input_data);
    assign temp_2 = ($unsigned((($signed(($unsigned(($signed(($signed(($unsigned(input_data) + (~input_data))) + temp_1[16:6])) | input_data)) + temp_1)) - (~input_data)) - temp_1)) | (~temp_0));
    assign temp_3 = ($signed(($signed(($signed(($signed(input_data) & input_data)) & temp_2[7:2])) & input_data)) & 32'd3361672518);
    assign temp_4 = (($signed((($signed(($signed((($unsigned(($signed(temp_0) | temp_2)) | input_data) + temp_3)) | input_data)) * temp_2) * (~temp_0))) - input_data) ^ input_data);
    assign temp_5 = $unsigned((($signed(($signed((($signed(temp_0) ^ temp_3) & temp_1)) & input_data)) * temp_3) + temp_2));
    logic [32:0] expr_331422;
    assign expr_331422 = ($unsigned((($unsigned(temp_4) + temp_2) ^ temp_5)) ^ temp_5);
    assign temp_6 = expr_331422[24:0];
    assign temp_7 = ($unsigned((($signed(($unsigned(($signed(($unsigned(((temp_1 + input_data) & input_data)) & input_data)) | temp_5)) & temp_1)) ^ input_data) - input_data)) + input_data);
    assign temp_8 = ($signed(($unsigned(($unsigned(($signed((temp_1 | temp_2)) + temp_6)) + temp_1)) - input_data)) & input_data);
    assign temp_9 = ((($signed(($unsigned(($unsigned(($unsigned((($signed(temp_3) - temp_0) - temp_4)) - temp_7)) + input_data)) ^ temp_8)) * temp_7) | temp_6) ^ input_data);
    assign temp_10 = ((((temp_3[31:13] | temp_6) ^ temp_3) ^ temp_6) | temp_4);
    assign temp_11 = {24'b0, (($signed(($signed(($unsigned(($signed((($unsigned((temp_6[24:15] + temp_2)) & temp_3) ^ temp_8)) <= temp_9)) >= temp_3)) >= temp_6)) >= temp_2) != temp_4)};
    logic [38:0] expr_286880;
    assign expr_286880 = $unsigned(((($signed((($unsigned(($signed((temp_9 ^ temp_11)) ^ temp_1)) - input_data) ^ (~temp_7))) + temp_5) ^ (~temp_0)) & (~temp_1)));
    assign temp_12 = expr_286880[27:0];
    assign temp_13 = (((((($unsigned(temp_11) & temp_6) * temp_9) << temp_11) - temp_1) + (~temp_8)) + temp_2);
    assign temp_14 = (($signed(((($unsigned(temp_11) | temp_12) & temp_5) * temp_7)) + temp_13) << temp_9);

    assign output_data = ($unsigned(((($unsigned((($unsigned(($signed(($unsigned(temp_2) * temp_9)) & (~temp_13))) & temp_9) ^ temp_5)) - temp_0) & temp_11) ^ temp_1[16:3])) - temp_10);

endmodule