module top (
    input [5:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;

    assign temp_0 = ((((((input_data | input_data) + input_data) + input_data) ^ input_data) + input_data) | input_data);
    assign temp_1 = $unsigned(temp_0);
    assign temp_2 = $signed(((((((temp_0 - temp_1) ^ temp_0) - temp_0) - temp_1[8:2]) + temp_1) | temp_0));
    assign temp_3 = $signed((((temp_2 & temp_0) & temp_2) + temp_1));
    assign temp_4 = temp_0 ? ((((input_data <= temp_3) - temp_3) ^ input_data) ^ input_data) : ((temp_2 * temp_1) + temp_2);
    assign temp_5 = ((temp_2 | temp_1) & input_data);
    assign temp_6 = (temp_0 | (~16'd8647));
    logic [26:0] expr_969964;
    assign expr_969964 = ((temp_0 * temp_2) & temp_2);
    assign temp_7 = expr_969964[13:0];
    assign temp_8 = (((((temp_2 * temp_3) - input_data) - temp_0) & temp_5) | temp_4);
    assign temp_9 = $signed(((((temp_2 + temp_0[12:0]) & temp_2[12:3]) & temp_1) * input_data[3:2]));
    assign temp_10 = $unsigned(((temp_0 ^ temp_5) & temp_4));
    assign temp_11 = (((temp_7 - temp_1) & temp_8) + temp_10);
    assign temp_12 = temp_0;
    assign temp_13 = $unsigned(temp_1);
    assign temp_14 = $unsigned((((temp_6 - temp_10) | (~temp_0)) + temp_5));

    assign output_data = $unsigned((temp_3 ^ temp_13));

endmodule