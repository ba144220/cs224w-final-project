module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;

    assign temp_0 = $signed(input_data);
    assign temp_1 = (temp_0 + input_data);
    assign temp_2 = {24'b0, temp_0};
    assign temp_3 = (temp_0 & input_data);
    assign temp_4 = (temp_1 | temp_0);
    logic [5:0] expr_46973;
    assign expr_46973 = (temp_4[5:5] - input_data[5:1]);
    assign temp_5 = expr_46973[4:0];
    assign temp_6 = $signed((temp_0 - temp_0));
    assign temp_7 = input_data;
    assign temp_8 = $signed(temp_6);
    assign temp_9 = temp_5;
    assign temp_10 = ((temp_3 - temp_7) ^ temp_4);
    logic [26:0] expr_918996;
    assign expr_918996 = $unsigned((input_data - temp_7));
    assign temp_11 = expr_918996[23:0];
    assign temp_12 = (temp_8 - temp_5);
    assign temp_13 = {10'b0, temp_2[30:29]};
    assign temp_14 = temp_12;
    assign temp_15 = temp_8;

    assign output_data = $unsigned(temp_15);

endmodule