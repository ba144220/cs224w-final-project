module top (
    input [2:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;
    logic [25:0] temp_16;
    logic [5:0] temp_17;
    logic [31:0] temp_18;

    assign temp_0 = input_data;
    assign temp_1 = input_data[1:1] ? $unsigned(temp_0) : ($signed(((($unsigned(temp_0) * temp_0[20:0]) ^ input_data) * temp_0)) * temp_0);
    assign temp_2 = $signed(input_data);
    assign temp_3 = (temp_2 | temp_2[2:0]);
    assign temp_4 = ((($unsigned(temp_0) ^ temp_2) | temp_1) | temp_3);
    assign temp_5 = temp_2[12:1];
    assign temp_6 = ((((temp_3 ^ temp_4) & temp_5) * input_data) & input_data);
    assign temp_7 = $signed(input_data);
    assign temp_8 = ((((temp_5 | temp_1[8:5]) | temp_4) ^ temp_5) - temp_3);
    assign temp_9 = temp_4[4:0];
    assign temp_10 = $unsigned(((((temp_1[8:2] - temp_5[8:4]) * temp_5[8:2]) & temp_4) | temp_4));
    assign temp_11 = ((temp_1 - input_data) - temp_0);
    assign temp_12 = ((temp_5 - temp_10) ^ input_data);
    assign temp_13 = $signed(((($unsigned(temp_5) & temp_9) - temp_6) | temp_9));
    assign temp_14 = (((temp_12 ^ temp_2) - temp_7) + temp_11);
    assign temp_15 = temp_9;
    assign temp_16 = $unsigned(((((temp_5 + temp_9) - temp_0[23:0]) + input_data) + temp_6));
    assign temp_17 = $unsigned((($unsigned(($signed(temp_13) - temp_11)) + temp_15) * temp_0));
    assign temp_18 = $unsigned((((temp_2 | temp_14) & temp_16) - temp_6));

    assign output_data = (((temp_12 + temp_12) + temp_15) + temp_0);

endmodule