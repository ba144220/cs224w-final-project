module top (
    input [3:0] input_data,
    output [36:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;

    assign temp_0 = 1'd1 ? {1'b0, input_data} : input_data;
    assign temp_1 = ($signed(($unsigned((temp_0 + (~temp_0))) * (~input_data))) * input_data);
    assign temp_2 = (($unsigned(temp_0) > input_data) < input_data);
    assign temp_3 = (($signed(temp_1) ^ temp_2) & input_data);
    assign temp_4 = temp_2[7:2] ? $signed(($signed(temp_2) + temp_0)) : $signed((($signed(temp_2) & temp_2) | (~input_data)));
    assign temp_5 = $unsigned(($unsigned((($unsigned(input_data) - (~temp_0)) * temp_1)) * temp_3));
    assign temp_6 = temp_5;
    assign temp_7 = ($unsigned((($unsigned(temp_2[2:0]) ^ temp_4) <= temp_6)) != temp_1);

    assign output_data = ((temp_7 + temp_5) - (~temp_5));

endmodule