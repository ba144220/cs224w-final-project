module top (
    input [4:0] input_data,
    output [36:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;
    logic [0:0] temp_13;

    assign temp_0 = $signed(($unsigned(($unsigned(($unsigned((input_data + 5'd0)) - input_data)) | input_data)) + input_data));
    assign temp_1 = ($signed(($signed(($signed(($signed(($unsigned(($unsigned(temp_0) | temp_0)) ^ input_data)) | input_data)) | temp_0)) | temp_0)) ^ temp_0);
    assign temp_2 = (($signed((($signed(($unsigned(((temp_1[16:8] ^ temp_0) * temp_0[4:1])) * temp_0)) * temp_1) & input_data)) - (~input_data)) - temp_1);
    logic [33:0] expr_174643;
    assign expr_174643 = $signed((($signed(($signed(($signed(($signed(($unsigned(temp_1) - input_data)) & temp_0[1:0])) & temp_2[7:2])) & temp_1)) & 32'd3361672518) & input_data));
    assign temp_3 = expr_174643[31:0];
    logic [34:0] expr_702977;
    assign expr_702977 = ($signed(($unsigned(($signed(temp_2) * (~temp_3))) - input_data)) * temp_2);
    assign temp_4 = expr_702977[28:0];
    assign temp_5 = temp_0 ? ($unsigned(($unsigned(($signed(((($signed(($signed((($unsigned(temp_1) << input_data) & temp_0[3:0])) << temp_0)) >> temp_2) - input_data) | temp_1)) ^ temp_4)) - temp_0[4:1])) * temp_2) : ($unsigned(temp_1) ^ temp_2);
    assign temp_6 = $signed(($unsigned(($unsigned((($signed(($unsigned(($signed(($unsigned((temp_2 & input_data)) & input_data)) | temp_5)) & temp_1)) ^ input_data) - temp_2)) ^ temp_0)) - temp_5));
    assign temp_7 = ($unsigned((($signed(($unsigned(($unsigned((temp_4 & temp_5)) + temp_0)) - input_data)) & (~input_data)) & input_data)) * (~temp_5));
    logic [30:0] expr_524677;
    assign expr_524677 = ($unsigned(($unsigned(temp_4) - temp_7)) + 7'd3);
    assign temp_8 = expr_524677[6:0];
    assign temp_9 = ($unsigned(($unsigned(((temp_5[15:0] ^ temp_4) + temp_6)) ^ temp_8)) ^ input_data);
    assign temp_10 = ($signed(($signed(($unsigned(($signed((($signed(input_data[1:0]) & input_data[3:2]) ^ temp_6)) | temp_4)) * (~temp_7))) + temp_0)) * temp_3);
    assign temp_11 = $signed(($signed(($unsigned(($signed((($signed(($signed(($unsigned((temp_8 - temp_6)) - temp_9)) * temp_3)) & (~temp_2)) ^ temp_4)) * (~temp_3))) | temp_3)) & temp_4));
    assign temp_12 = ($signed(($signed((((($signed(($signed(temp_4) - 28'd257911948)) - temp_10) + temp_4) + temp_8[6:3]) - temp_10)) & temp_10)) | temp_6);
    logic [37:0] expr_684274;
    assign expr_684274 = (($unsigned(((((temp_9 | temp_1) + (~temp_8)) + temp_2) | (~temp_12))) | (~temp_2)) & temp_3);
    assign temp_13 = expr_684274[0:0];

    assign output_data = $signed((($unsigned(($signed(($signed(((($unsigned(($signed(temp_13) + temp_13)) & temp_5) & temp_4) + temp_8)) | temp_1)) & (~temp_13))) & temp_9) ^ temp_5));

endmodule