module top (
    input [4:0] input_data,
    output [9:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;
    logic [26:0] temp_10;
    logic [4:0] temp_11;
    logic [15:0] temp_12;
    logic [5:0] temp_13;
    logic [27:0] temp_14;
    logic [3:0] temp_15;
    logic [7:0] temp_16;
    logic [14:0] temp_17;

    assign temp_0 = ($unsigned(($signed(input_data) + (~input_data))) * input_data);
    assign temp_1 = ($signed(($unsigned(input_data[4:1]) * temp_0)) ^ input_data[3:0]);
    assign temp_2 = input_data[4:4] ? ($unsigned(input_data) + input_data) : ($unsigned(temp_1) & temp_1[1:0]);
    assign temp_3 = ($signed(input_data) * input_data);
    assign temp_4 = ($unsigned(input_data) - input_data);
    assign temp_5 = $unsigned(($signed(temp_0) + temp_0[19:0]));
    assign temp_6 = (temp_0 & temp_2[1:0]);
    assign temp_7 = temp_4;
    assign temp_8 = input_data[1:1] ? (input_data | input_data) : input_data;
    assign temp_9 = $unsigned(($unsigned(input_data) + temp_3));
    assign temp_10 = (($signed(temp_3) ^ temp_6) + temp_7);
    assign temp_11 = temp_1;
    assign temp_12 = temp_9;
    assign temp_13 = (temp_8[2:0] | (~temp_7));
    assign temp_14 = temp_10 ? temp_0 : temp_8;
    assign temp_15 = input_data[3:0];
    assign temp_16 = temp_13[3:0];
    assign temp_17 = ($unsigned((temp_4 + (~temp_15[3:0]))) & (~temp_12));

    assign output_data = temp_10 ? {7'b0, temp_7} : temp_13;

endmodule