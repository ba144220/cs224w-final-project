module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;

    assign temp_0 = ((input_data | input_data) * input_data);
    assign temp_1 = temp_0 ? ($signed(((((((($unsigned(temp_0) * input_data) & temp_0) * temp_0) ^ temp_0) | temp_0) | temp_0) | input_data)) - 24'd1641151) : $signed((($unsigned(($unsigned(($signed(input_data) + (~temp_0))) + temp_0)) + input_data) ^ temp_0));
    assign temp_2 = ((temp_1 - temp_1) * temp_1);
    assign temp_3 = temp_0 ? temp_1[8:0] : (($unsigned(((($signed(temp_0) - temp_2[2:0]) - temp_2) - temp_1)) | (~temp_0)) * (~temp_1));
    assign temp_4 = $unsigned((($signed(($signed(($signed((($unsigned(($signed(temp_0[1:0]) ^ temp_0)) * temp_3) < input_data)) + temp_3)) > temp_3)) | temp_0) * temp_0));
    assign temp_5 = ((($signed(($signed(($signed(temp_4) & temp_4)) - (~temp_2))) | temp_1) & temp_3) + temp_1);
    assign temp_6 = ((($signed((($unsigned(((($unsigned(temp_0[2:0]) ^ temp_3) - (~temp_4)) ^ temp_2)) + temp_3) * temp_4)) & temp_5) & (~temp_1[18:0])) + temp_3);

    assign output_data = ((($unsigned((temp_2 | temp_5)) & (~temp_3)) + (~temp_1)) - temp_0);

endmodule