module top (
    input [2:0] input_data,
    output [18:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;
    logic [0:0] temp_13;
    logic [28:0] temp_14;
    logic [17:0] temp_15;

    assign temp_0 = {1'b0, $signed((input_data + input_data))};
    assign temp_1 = $unsigned((((temp_0 + (~temp_0)) * input_data) - (~temp_0)));
    assign temp_2 = ((temp_0 & input_data) | input_data);
    assign temp_3 = (input_data ^ temp_2[7:0]);
    assign temp_4 = $unsigned((input_data << temp_2));
    assign temp_5 = (input_data + input_data);
    assign temp_6 = (temp_4 | temp_2);
    assign temp_7 = (input_data - temp_1);
    assign temp_8 = (((temp_5 ^ temp_3) * temp_6) | input_data);
    assign temp_9 = (((temp_6 << temp_7) * temp_5) | temp_6);
    assign temp_10 = input_data[2:1];
    assign temp_11 = ((temp_9 >> temp_8) * (~temp_5));
    logic [32:0] expr_955005;
    assign expr_955005 = (($signed(input_data) + temp_4) + temp_9);
    assign temp_12 = expr_955005[27:0];
    assign temp_13 = ((temp_3 + temp_4) + temp_9);
    assign temp_14 = $unsigned(((temp_3 + input_data) * temp_2));
    assign temp_15 = $unsigned((temp_4 + temp_0));

    assign output_data = (temp_4 + temp_9);

endmodule