module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;

    assign temp_0 = ($unsigned((input_data + input_data)) * input_data);
    assign temp_1 = input_data;
    assign temp_2 = ((((temp_1 + temp_1) * temp_0[2:0]) - temp_1) ^ (~temp_0));
    assign temp_3 = ((temp_1 ^ temp_2) * temp_1);
    logic [31:0] expr_441682;
    assign expr_441682 = $signed(((temp_1[25:24] - temp_1) + temp_2));
    assign temp_4 = expr_441682[5:0];
    assign temp_5 = $unsigned((((((temp_0[3:0] - temp_1) * temp_4) ^ temp_3) - temp_3) ^ temp_2));
    assign temp_6 = ($unsigned((((temp_0 & temp_5) - temp_2) | temp_1)) & input_data[1:0]);
    assign temp_7 = temp_6 ? (($signed(temp_4) * temp_6) * temp_3) : $unsigned(((($signed(temp_6) * temp_2) + temp_3) & (~temp_2)));
    assign temp_8 = ((($unsigned(($unsigned(temp_7) | temp_5)) * temp_5) * temp_5) + temp_1);
    assign temp_9 = $unsigned(temp_3);
    assign temp_10 = ($unsigned(((temp_5 & temp_6) | temp_2)) & temp_9[3:0]);

    assign output_data = temp_10;

endmodule