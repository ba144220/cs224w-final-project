module top (
    input [5:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;

    assign temp_0 = input_data;
    assign temp_1 = (temp_0 + input_data);
    assign temp_2 = input_data;
    assign temp_3 = (temp_2 ^ temp_2);
    assign temp_4 = ((temp_0 + temp_3) + (~temp_0));
    assign temp_5 = $unsigned((temp_3 * input_data));
    assign temp_6 = {5'b0, ((temp_3 | temp_2[8:0]) + input_data)};
    assign temp_7 = $signed((temp_0 - temp_4));
    assign temp_8 = temp_0;
    assign temp_9 = (($signed(temp_3) | temp_0) & temp_4);
    assign temp_10 = (temp_3 | temp_4);
    assign temp_11 = ((temp_7 + temp_1) | temp_4);
    assign temp_12 = temp_3;
    logic [29:0] expr_200533;
    assign expr_200533 = $unsigned(temp_12);
    assign temp_13 = expr_200533[24:0];

    assign output_data = $unsigned(temp_10);

endmodule