module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;

    assign temp_0 = $signed(input_data);
    assign temp_1 = $unsigned(($signed(input_data) & input_data));
    assign temp_2 = ($unsigned(temp_0) * (~input_data));
    assign temp_3 = temp_2;
    assign temp_4 = ($signed(($signed(temp_1[25:12]) ^ temp_2)) ^ temp_0);
    assign temp_5 = temp_1 ? $unsigned((temp_1[25:24] - temp_1)) : $signed(($signed(temp_3[9:7]) & temp_3));
    assign temp_6 = temp_2 ? $unsigned((input_data[1:0] & temp_3)) : $unsigned(((temp_5 & input_data[2:1]) + (~temp_4)));
    assign temp_7 = $unsigned((26'd15554488 << input_data));
    assign temp_8 = $unsigned((($unsigned(temp_0) + temp_4[5:3]) * input_data));
    assign temp_9 = (temp_5 != temp_1);
    assign temp_10 = $signed(($unsigned(temp_7) + temp_0[6:1]));
    assign temp_11 = temp_9;
    assign temp_12 = $signed(($unsigned((temp_2 ^ temp_6)) * temp_5));
    assign temp_13 = $unsigned(((temp_12 - (~temp_9)) - temp_7));
    assign temp_14 = $unsigned(($signed(temp_5) & temp_6));

    assign output_data = (temp_0[6:6] * temp_9);

endmodule