module top (
    input [2:0] input_data,
    output [7:0] output_data
);

    logic [16:0] temp_0;
    logic [2:0] temp_1;
    logic [0:0] temp_2;
    logic [9:0] temp_3;
    logic [30:0] temp_4;
    logic [23:0] temp_5;
    logic [20:0] temp_6;
    logic [1:0] temp_7;
    logic [17:0] temp_8;
    logic [31:0] temp_9;
    logic [12:0] temp_10;
    logic [26:0] temp_11;
    logic [6:0] temp_12;
    logic [12:0] temp_13;
    logic [16:0] temp_14;

    assign temp_0 = $signed(($unsigned(($unsigned(($signed(($signed(($unsigned(((($signed((input_data * input_data)) - input_data) ^ input_data) | input_data)) & input_data)) + input_data)) - input_data)) | input_data)) ^ input_data));
    assign temp_1 = temp_0 ? ($unsigned(temp_0) ^ temp_0) : ((((((((temp_0 & temp_0) ^ input_data) & temp_0) * temp_0) ^ temp_0) - input_data) | temp_0) - (~temp_0[4:0]));
    assign temp_2 = temp_0 ? ((input_data[1:1] & temp_0) & temp_1) : $signed(temp_1);
    assign temp_3 = ((((((($unsigned(($signed(temp_0[7:0]) ^ temp_0)) ^ temp_0) ^ temp_2) ^ input_data) | temp_2) + temp_2) ^ temp_2) + temp_0);
    assign temp_4 = temp_3 ? ((($signed(($unsigned(temp_0) - input_data)) == input_data) == temp_1[2:2]) >= (~temp_2)) : (($unsigned((((($signed(temp_0[3:0]) & temp_2) - temp_3) * temp_2) | temp_0)) | temp_3) + temp_2);
    assign temp_5 = ((((((24'd4223166 - temp_0) * input_data) + temp_0) | temp_0) * temp_1) ^ input_data);
    assign temp_6 = ($signed(($unsigned((($unsigned(temp_5[21:0]) & temp_0) * temp_1)) | input_data)) - temp_3);
    assign temp_7 = ((($unsigned(($unsigned(($signed((($signed((temp_2 ^ (~temp_4))) & temp_2) - temp_2)) ^ temp_0)) ^ temp_3)) + (~temp_4)) ^ temp_6) & temp_0);
    assign temp_8 = ($unsigned(((($unsigned(($signed(($signed((($unsigned(temp_6) | temp_1) != temp_1)) & temp_0)) == temp_0)) > temp_4) >= temp_6) >= temp_2)) >= temp_4);
    assign temp_9 = (temp_7 & (~temp_5));
    assign temp_10 = (($unsigned(((((($unsigned(temp_5) & temp_1) & temp_0) * (~input_data)) | temp_0) | (~temp_4))) * temp_2) + temp_7);
    assign temp_11 = $signed((temp_4 * temp_10));
    assign temp_12 = temp_10;
    assign temp_13 = (temp_10 + (~temp_3));
    assign temp_14 = (((temp_12 & temp_9) - (~temp_13)) & temp_4);

    assign output_data = (($unsigned((((temp_12 | temp_4) + (~temp_2)) - (~temp_8))) & temp_1) * (~temp_12));

endmodule