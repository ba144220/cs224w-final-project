module top (
    input [3:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;

    assign temp_0 = (($unsigned((25'd27357858 & input_data)) + (~input_data)) + input_data);
    assign temp_1 = temp_0 ? (($signed(($unsigned((temp_0 - input_data)) & temp_0)) | input_data) * temp_0) : ($unsigned(($unsigned((($signed((input_data + input_data)) * (~temp_0[24:3])) - input_data)) * -9'd36)) | (~temp_0[16:0]));
    assign temp_2 = (($unsigned(($signed(($unsigned(temp_0[20:0]) - temp_1)) ^ temp_0)) - temp_0[24:0]) ^ temp_1);
    assign temp_3 = ((3'd1 ^ temp_1) * input_data[3:1]);
    assign temp_4 = input_data;
    assign temp_5 = $unsigned((($unsigned(($unsigned((($unsigned(temp_4) - temp_4[5:2]) & input_data)) | temp_3)) - input_data) & temp_1));
    assign temp_6 = temp_5 ? 16'd11004 : ((($unsigned(($signed((temp_1 * (~temp_5))) ^ temp_3)) + (~temp_0[24:24])) ^ temp_1) & temp_5);
    assign temp_7 = (($unsigned((temp_4 & temp_5)) * input_data) - input_data);
    assign temp_8 = (((temp_5 & temp_2[12:3]) & temp_1) * input_data);
    assign temp_9 = ((temp_0 ^ input_data[1:0]) & temp_8[25:9]);
    assign temp_10 = ((temp_1 * temp_1) & (~temp_8[25:5]));
    assign temp_11 = (temp_3[2:2] ^ temp_5);
    assign temp_12 = temp_5[8:4] ? temp_3 : temp_11;
    assign temp_13 = temp_0;
    assign temp_14 = temp_8[25:7];

    assign output_data = temp_13;

endmodule