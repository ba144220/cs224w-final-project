module top (
    input [2:0] input_data,
    output [4:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;

    assign temp_0 = input_data;
    assign temp_1 = ((($signed((($signed(temp_0) - input_data) | input_data)) > temp_0) <= temp_0[6:6]) & temp_0);
    assign temp_2 = temp_0;
    assign temp_3 = (input_data * temp_0);
    assign temp_4 = (((((((temp_1[25:2] & temp_2) - temp_0[6:6]) | temp_1[25:17]) ^ input_data) - temp_1) + temp_1) * temp_2);
    assign temp_5 = ((((($unsigned(((input_data * temp_3) ^ input_data)) + input_data) * temp_0) & input_data) | input_data) - temp_4);
    assign temp_6 = (((((((($unsigned((temp_1[25:17] + temp_2[30:18])) * temp_3) * temp_3) - temp_3) - temp_2) ^ temp_5) & temp_4) ^ temp_0) | temp_4);
    assign temp_7 = ($signed(($signed(temp_4) * temp_6)) - temp_2);
    assign temp_8 = (temp_1 + temp_7);
    assign temp_9 = (((((((((temp_5 ^ temp_7) * temp_0) * temp_6[1:1]) ^ input_data) & temp_7) * temp_0) | temp_8) + temp_0) - temp_6);
    assign temp_10 = ((((((($signed((temp_8[18:9] | temp_4)) + temp_0) + temp_8[18:0]) ^ temp_6) & temp_5) + temp_3) & temp_5[4:2]) ^ 15'd31204);
    assign temp_11 = ((((((((temp_10 - temp_1) + temp_9) + temp_2) * (~temp_10[14:7])) | temp_4) * temp_0) & input_data) * temp_1[9:0]);
    assign temp_12 = ($unsigned((($signed(((((($signed(((((temp_4 >> temp_10) & temp_1) * temp_1) * temp_4[3:0])) ^ input_data) + (~temp_4)) & temp_6) << temp_0) & input_data)) & temp_5) ^ input_data)) << temp_6);
    assign temp_13 = ((($unsigned(temp_1) | temp_9) - temp_2[30:20]) * temp_5);
    assign temp_14 = (((((temp_9 >> temp_1) * temp_0) + temp_9) | (~temp_7)) * temp_6);
    assign temp_15 = (($signed((((($unsigned((((((($signed(temp_13) - temp_14[6:1]) | temp_1) | temp_0[6:4]) | temp_5[4:1]) | temp_2) | temp_12)) & temp_7) * temp_10) - temp_5) | temp_5[4:1])) * temp_3[9:5]) + temp_10);

    assign output_data = $unsigned((((((((((((temp_10[14:1] & temp_0[6:6]) * temp_10) + temp_12) ^ temp_2[30:13]) + temp_9[3:2]) & temp_10) ^ temp_3) + temp_15) | (~temp_5)) ^ temp_7) & temp_14));

endmodule