module top (
    input [11:0] input_data,
    output [2:0] output_data
);

    logic [31:0] temp_0;
    logic [16:0] temp_1;
    logic [2:0] temp_2;
    logic [0:0] temp_3;
    logic [9:0] temp_4;
    logic [30:0] temp_5;
    logic [23:0] temp_6;
    logic [20:0] temp_7;
    logic [1:0] temp_8;
    logic [17:0] temp_9;
    logic [31:0] temp_10;
    logic [12:0] temp_11;
    logic [26:0] temp_12;

    assign temp_0 = $unsigned((input_data ^ input_data));
    assign temp_1 = ($unsigned(input_data) | input_data);
    assign temp_2 = $unsigned(temp_1[16:7]);
    logic [22:0] expr_395814;
    assign expr_395814 = ($signed(($signed((($unsigned((($signed(($unsigned(input_data[8:8]) + temp_0[11:0])) * temp_1) & temp_1)) & temp_1) + temp_2)) + temp_1)) * input_data[6:6]);
    assign temp_3 = expr_395814[0:0];
    assign temp_4 = (($unsigned(($signed(($signed(($unsigned(($unsigned((input_data[10:1] ^ temp_2)) * temp_3)) * temp_3)) & (~input_data[11:2]))) * input_data[9:0])) + input_data[10:1]) ^ temp_0[21:0]);
    assign temp_5 = ($signed((input_data & temp_3)) * temp_0[28:0]);
    assign temp_6 = (($unsigned((temp_0 + temp_5)) + temp_5[18:0]) - temp_4);
    assign temp_7 = ($unsigned(($unsigned((temp_1 * input_data)) - temp_6)) ^ temp_1);
    assign temp_8 = $signed(temp_1);
    assign temp_9 = ($signed(($unsigned((($signed(temp_0[22:0]) > temp_1) != temp_4)) <= temp_3)) != temp_5[30:20]);
    logic [34:0] expr_437877;
    assign expr_437877 = ($unsigned(($unsigned((($unsigned(($signed(temp_2[2:0]) + temp_7[20:19])) | temp_6) * temp_0)) + temp_1[13:0])) ^ temp_7);
    assign temp_10 = expr_437877[31:0];
    assign temp_11 = ($signed(($signed(temp_3) + temp_9)) - temp_0);
    assign temp_12 = ($unsigned(temp_9) | temp_11);

    assign output_data = ($signed(($unsigned(($unsigned(temp_10[16:0]) ^ temp_7)) * temp_11[6:0])) + temp_0[31:21]);

endmodule