module top (
    input [3:0] input_data,
    output [34:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;

    assign temp_0 = ((input_data - (~input_data)) * input_data);
    assign temp_1 = ((temp_0 ^ input_data) & temp_0);
    assign temp_2 = ((((((((temp_0 * temp_0) + (~temp_0)) | temp_0) * temp_0[8:1]) * temp_0) - input_data) | temp_0) ^ temp_1);
    assign temp_3 = $unsigned(((((((temp_2 * (~temp_1[23:2])) * temp_1) * input_data) | temp_0) - temp_2[30:11]) - temp_0));
    assign temp_4 = (((((temp_2 + input_data[1:1]) * temp_3) - (~temp_3)) & input_data[2:2]) + (~input_data[0:0]));
    assign temp_5 = ((((((temp_1 + (~temp_3)) | temp_0) - (~temp_2)) ^ temp_3) & (~temp_2[30:2])) + temp_0[8:8]);
    assign temp_6 = (((((temp_1 & temp_4) & temp_0) ^ temp_5[30:7]) + temp_1) | temp_2);
    assign temp_7 = (temp_4 - temp_0);
    assign temp_8 = $unsigned(temp_4);
    assign temp_9 = $unsigned((temp_8 + temp_2));
    assign temp_10 = $unsigned((temp_2 | (~temp_8[12:7])));
    assign temp_11 = (((((((temp_3 - temp_8) | temp_4) - temp_5) ^ temp_9) + temp_1) & temp_3) * temp_3[4:1]);
    assign temp_12 = (((((((((((temp_4 ^ (~temp_0)) ^ temp_7) ^ temp_7) * temp_5) * temp_5) * temp_4) ^ temp_5) - temp_10) & temp_2[30:6]) ^ (~temp_1)) | temp_11);

    assign output_data = (temp_10 != temp_1);

endmodule