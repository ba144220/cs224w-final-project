module top (
    input [2:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;

    assign temp_0 = ($signed(($unsigned(($signed(($unsigned(input_data) * (~input_data))) ^ input_data)) ^ input_data)) | input_data);
    assign temp_1 = (($signed((($unsigned(input_data) < (~temp_0)) + temp_0)) == temp_0) >= temp_0[6:1]);
    assign temp_2 = ($signed(($signed(temp_0) ^ temp_1[10:0])) | temp_0);
    assign temp_3 = input_data;
    assign temp_4 = (temp_1 >= temp_0);
    assign temp_5 = (($unsigned((((($unsigned(temp_3) + temp_2) + input_data) ^ temp_0[6:2]) - temp_3)) ^ temp_2) ^ temp_0);
    assign temp_6 = ($unsigned(($unsigned(($signed((($signed(((temp_1 - temp_2) | temp_1)) & temp_3[1:0]) * temp_1[3:0])) + temp_2[30:18])) & temp_3)) * temp_3);
    assign temp_7 = ($signed(temp_1) * temp_0[6:3]);

    assign output_data = (($unsigned(($unsigned(($unsigned(($unsigned((temp_2 ^ temp_0)) | temp_4)) * temp_5)) | temp_2)) + temp_1) * (~temp_0));

endmodule