module top (
    input [2:0] input_data,
    output [36:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;
    logic [0:0] temp_13;
    logic [28:0] temp_14;
    logic [17:0] temp_15;
    logic [14:0] temp_16;
    logic [6:0] temp_17;
    logic [20:0] temp_18;

    assign temp_0 = 1'd1 ? ($signed((($signed(input_data) & input_data) * input_data)) ^ input_data) : $unsigned(((($unsigned(($unsigned(($unsigned((input_data | input_data)) | input_data)) - (~input_data))) - input_data) * (~input_data)) - input_data));
    assign temp_1 = $unsigned(($unsigned(($signed(($signed(($unsigned((($unsigned(($signed(input_data) ^ temp_0)) | temp_0) | (~temp_0))) + (~input_data))) + (~temp_0[4:2]))) | input_data)) + temp_0));
    assign temp_2 = temp_0[2:0] ? $signed(($signed(($unsigned(($unsigned(($unsigned(($unsigned(((temp_0 ^ temp_0[4:3]) ^ temp_0)) * input_data)) | input_data)) ^ 8'd50)) - temp_1)) + temp_1)) : $signed(((($unsigned(($signed(((($unsigned(($signed(temp_0) | temp_1)) | (~input_data)) + temp_1) | temp_1)) * input_data)) * temp_0[4:1]) - temp_0) & input_data));
    assign temp_3 = input_data[2:2] ? ($signed(($unsigned(($unsigned((($signed((($signed(($signed((temp_0 & temp_0)) & (~input_data))) * temp_1) + temp_1)) + (~temp_2[7:2])) | input_data)) * temp_0)) - input_data)) | temp_0) : $signed(($signed(($unsigned((temp_2 + input_data)) | temp_1)) | temp_2));
    assign temp_4 = $signed(input_data);
    assign temp_5 = ((($signed(((($unsigned(input_data) + input_data) * temp_2) | (~temp_0))) * temp_4) & (~temp_1)) * temp_2[7:2]);
    assign temp_6 = input_data[1:1] ? (($unsigned((($unsigned((($signed(temp_4) + temp_4[28:10]) - temp_4[21:0])) * temp_2) & input_data)) + input_data) + temp_5[10:0]) : ($signed((($unsigned(((((($unsigned(temp_5) + temp_5) & temp_3) ^ input_data) | temp_5) ^ temp_2)) * input_data) ^ temp_0)) * input_data);
    assign temp_7 = $signed(($unsigned((((temp_4 + (~temp_5)) + temp_5) * temp_0)) | input_data));
    assign temp_8 = ((($signed(temp_0) & temp_6) | (~temp_2)) - input_data);
    assign temp_9 = ($unsigned(input_data) + 32'd2934748484);
    assign temp_10 = $signed(($unsigned(((($unsigned(temp_6) * input_data[2:1]) != (~temp_7)) + input_data[2:1])) & (~temp_2[7:4])));
    assign temp_11 = input_data;
    assign temp_12 = $signed(($unsigned(($unsigned((((($signed(($unsigned(temp_3) ^ temp_4)) * temp_11) - temp_8) ^ (~input_data)) - temp_0[1:0])) | temp_5[18:0])) ^ (~input_data)));
    assign temp_13 = ((temp_10 - temp_3) | temp_2);
    assign temp_14 = ($unsigned((($unsigned(($signed(temp_5) | temp_4)) * temp_8) * temp_7)) & temp_1);
    assign temp_15 = ($unsigned(((((temp_6 * temp_2[3:0]) + temp_6) ^ temp_1[16:3]) - temp_2)) & temp_4);
    assign temp_16 = ($unsigned(((temp_8[6:5] & temp_15) & temp_14[10:0])) | temp_9);
    assign temp_17 = (($signed(((($signed((((temp_9 - temp_5[30:14]) * temp_9) + temp_12)) & temp_12[27:12]) * temp_4) | temp_13)) ^ temp_12[27:5]) + (~temp_15[17:6]));
    assign temp_18 = $signed(($unsigned((($unsigned((((($unsigned((temp_3 - (~temp_8))) & temp_2[7:4]) - temp_15) | temp_17) & temp_10[1:1])) | temp_14) & temp_4)) + temp_16));

    assign output_data = $unsigned(($unsigned(($unsigned(($unsigned(($signed((($signed(($signed(($unsigned((temp_18 + temp_16)) - temp_10)) - (~temp_2))) | temp_6) * temp_7)) * (~temp_8))) * temp_4[28:3])) - temp_8)) ^ temp_7));

endmodule