module top (
    input [4:0] input_data,
    output [36:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;

    assign temp_0 = input_data;
    assign temp_1 = temp_0 ? $unsigned(temp_0) : ($signed(input_data) - input_data);
    assign temp_2 = ($unsigned(($signed(input_data) | input_data)) ^ input_data);
    assign temp_3 = input_data;
    assign temp_4 = input_data;
    assign temp_5 = ($signed(input_data) | input_data);
    assign temp_6 = $unsigned(($unsigned(temp_4) - temp_4));
    assign temp_7 = temp_0 ? $signed(($signed(temp_0) - (~temp_5))) : {9'b0, input_data};
    assign temp_8 = temp_2 ? $unsigned(($unsigned(input_data) - (~temp_0))) : ($unsigned(input_data) << temp_2[7:0]);
    assign temp_9 = ($signed(($unsigned(temp_1) << (~temp_7[11:0]))) << 32'd3361672518);
    assign temp_10 = $signed(($unsigned(temp_8) + temp_2));
    assign temp_11 = $unsigned(($signed(($unsigned(temp_9[31:2]) & temp_2)) | temp_9[9:0]));
    assign temp_12 = temp_9[31:4] ? temp_2[2:0] : {21'b0, $signed(temp_8)};

    assign output_data = {8'b0, $signed(temp_4)};

endmodule