module top (
    input [5:0] input_data,
    output [18:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;

    assign temp_0 = (input_data ^ 9'd163);
    assign temp_1 = ((($signed(temp_0) & input_data) ^ input_data) | temp_0);
    assign temp_2 = {24'b0, ($signed(input_data) ^ input_data)};
    assign temp_3 = (((temp_1[23:20] + temp_2) + temp_0) | input_data[4:0]);
    assign temp_4 = (($signed(($unsigned(input_data[4:4]) + input_data[4:4])) * temp_2) + temp_1[21:0]);
    assign temp_5 = {6'b0, ((($unsigned(input_data) == temp_4) | temp_3) * temp_1)};
    assign temp_6 = (($unsigned(input_data) * (~input_data)) - temp_4);
    assign temp_7 = ((temp_5 & temp_3[4:4]) ^ temp_5);
    assign temp_8 = $unsigned(($signed(($unsigned(((((temp_0[4:0] & temp_0) + temp_6[4:0]) | temp_0) - (~temp_4))) ^ temp_6[9:0])) + temp_0));
    assign temp_9 = $signed((temp_4 * (~temp_2)));
    assign temp_10 = (((temp_0 ^ temp_6) + temp_3) | temp_4);
    assign temp_11 = temp_9;

    assign output_data = ((((temp_2 + temp_0) | temp_4) ^ (~temp_3)) * temp_9);

endmodule