module top (
    input [2:0] input_data,
    output [18:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;

    assign temp_0 = input_data;
    assign temp_1 = ((input_data != (~input_data)) ^ temp_0);
    assign temp_2 = $signed(((temp_1 * input_data) | input_data));
    assign temp_3 = (temp_0[7:0] & 5'd2);
    assign temp_4 = $signed(temp_0);
    assign temp_5 = $unsigned((input_data | temp_4));
    assign temp_6 = $unsigned((temp_0 * temp_4));
    assign temp_7 = $signed((temp_2 >= temp_1));
    assign temp_8 = temp_2 ? ($signed(temp_1[11:0]) * temp_3) : ($unsigned(temp_3) | temp_4);
    assign temp_9 = (temp_6[14:0] - temp_7);
    assign temp_10 = ($signed(($unsigned(temp_4) + temp_4)) - temp_6[16:4]);
    assign temp_11 = $unsigned((($unsigned(temp_8) * temp_1) - temp_0));

    assign output_data = $signed(temp_0);

endmodule