module top (
    input [4:0] input_data,
    output [4:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;
    logic [26:0] temp_10;
    logic [4:0] temp_11;

    assign temp_0 = {13'b0, $signed(($signed(((((($unsigned(($signed((input_data ^ input_data)) - (~input_data))) * input_data) + input_data) & input_data) & input_data) - input_data)) ^ input_data))};
    assign temp_1 = $unsigned(($signed((($signed(($signed(($signed(($unsigned(((temp_0 & (~temp_0)) ^ (~temp_0))) & temp_0)) & temp_0)) ^ (~temp_0))) ^ temp_0) | input_data[3:0])) ^ input_data[4:1]));
    assign temp_2 = input_data[4:4] ? ($signed((input_data | (~temp_1))) & input_data) : $signed((($signed(input_data) | temp_0) | temp_1));
    assign temp_3 = $unsigned((($signed((temp_0 - input_data)) * input_data) & temp_2));
    assign temp_4 = ((($signed(input_data) & temp_0) ^ (~temp_3)) + input_data);
    assign temp_5 = (((temp_4 * temp_2) <= temp_1) + input_data[3:0]);
    assign temp_6 = ($signed(($unsigned(((($signed((($unsigned((input_data * temp_0)) & temp_4) | input_data)) - input_data) & temp_5) ^ temp_1)) + temp_3)) & temp_1);
    assign temp_7 = ($signed((((input_data[2:0] - temp_0) | (~temp_4)) + temp_1)) | temp_6);
    assign temp_8 = temp_2;
    assign temp_9 = (((temp_5 + temp_8) + temp_6) * temp_3);
    assign temp_10 = temp_1 ? ((($signed((($unsigned((temp_8 & temp_0)) ^ input_data) * temp_6[5:0])) <= (~temp_1)) | temp_1) != (~temp_9)) : $unsigned(temp_6);
    assign temp_11 = $signed(temp_10);

    assign output_data = ($signed(($unsigned((($unsigned(($unsigned((temp_10[18:0] ^ temp_3)) | temp_8[5:0])) + temp_4) & temp_1)) ^ temp_3[2:0])) | temp_9[16:0]);

endmodule