module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;

    assign temp_0 = ((((input_data + input_data) & input_data) + 6'd46) - input_data);
    assign temp_1 = $unsigned(((temp_0 | temp_0) & input_data));
    assign temp_2 = (($unsigned(temp_1) | temp_0) + temp_0);
    assign temp_3 = {13'b0, (input_data ^ (~temp_0))};
    assign temp_4 = {10'b0, (temp_0 + temp_0)};
    assign temp_5 = $signed((((temp_1[22:0] * temp_0) & temp_2) & temp_4));
    assign temp_6 = temp_2[4:0];
    assign temp_7 = (($signed(temp_1[14:0]) - temp_5[2:0]) - temp_5);
    assign temp_8 = (((temp_6 - temp_7) | temp_5) & temp_0);
    assign temp_9 = temp_4 ? (((temp_7 + temp_1[11:0]) ^ temp_7) & temp_5) : ((temp_8 + temp_1[6:0]) & (~temp_1));

    assign output_data = ((temp_1 & temp_1) - temp_7);

endmodule