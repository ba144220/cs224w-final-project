module top (
    input [3:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;

    assign temp_0 = (((input_data ^ input_data) ^ 25'd4233809) + (~input_data));
    assign temp_1 = ((temp_0[19:0] & input_data) & temp_0);
    assign temp_2 = (((((temp_0 * temp_1[5:0]) & temp_1[1:0]) * temp_1) & (~temp_1)) + input_data);
    assign temp_3 = (((temp_2[5:0] ^ temp_1[8:0]) + input_data[2:0]) > temp_0);
    assign temp_4 = ((temp_3 & temp_1[2:0]) ^ temp_0);
    assign temp_5 = (((((((((temp_4[5:5] * input_data) | temp_2) * input_data) | input_data) ^ temp_2) & (~input_data)) ^ input_data) * temp_4) - input_data);
    assign temp_6 = (temp_4 - temp_1);
    assign temp_7 = ((((($unsigned(((((temp_6[15:0] + (~input_data)) - temp_4) + temp_0) & temp_5)) - temp_1[1:0]) - temp_2) ^ input_data) - temp_6) * temp_3);
    assign temp_8 = ((((((((input_data & temp_4) & temp_1[8:6]) & temp_2[12:3]) & temp_1) * input_data) - temp_7) * temp_0) + temp_3);
    assign temp_9 = temp_4 ? $signed(((((temp_1 * temp_1) & temp_8) + temp_4) - (~2'd1))) : $unsigned(((($unsigned((temp_5 & 2'd0)) << input_data[1:0]) ^ input_data[1:0]) & input_data[2:1]));
    assign temp_10 = ((((temp_3 ^ input_data) - temp_1) & input_data) & temp_8);
    assign temp_11 = (((temp_1 - temp_9[1:1]) + temp_10) & temp_3[1:0]);
    assign temp_12 = (((((((temp_0 | temp_3[2:2]) & temp_7) + temp_7) ^ temp_8) ^ temp_1) * temp_9) * temp_5[8:7]);
    assign temp_13 = (((((((temp_8[3:0] ^ temp_1) & (~temp_3)) * temp_8) * temp_1[8:0]) ^ temp_0) ^ temp_1) - temp_11);

    assign output_data = $signed(((((((((temp_5[3:0] <= temp_5) & temp_6) * temp_10[10:0]) - temp_7) < (~temp_5)) >= temp_10[18:0]) != temp_6[5:0]) + temp_10));

endmodule