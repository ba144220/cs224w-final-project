module top (
    input [3:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;
    logic [25:0] temp_16;
    logic [5:0] temp_17;

    assign temp_0 = (($unsigned((($signed(($unsigned(($unsigned(input_data) != 25'd4233809)) + input_data)) >= input_data) * input_data)) | input_data) != input_data);
    assign temp_1 = $unsigned(($signed(($signed(($unsigned(($signed(input_data) * temp_0)) ^ input_data)) + temp_0[24:13])) - temp_0[24:3]));
    assign temp_2 = ($signed(($signed(((temp_0[5:0] ^ (~temp_0)) >> temp_0)) * temp_1[8:4])) - temp_1);
    logic [10:0] expr_381784;
    assign expr_381784 = temp_2[10:0];
    assign temp_3 = expr_381784[2:0];
    assign temp_4 = ((($unsigned(($unsigned(input_data) <= temp_3)) != temp_3) != input_data) - temp_2);
    assign temp_5 = ($unsigned(($unsigned((($signed(input_data) ^ temp_3) * input_data)) | temp_3)) - input_data);
    assign temp_6 = $unsigned((($signed(($unsigned(temp_4) + temp_5)) ^ temp_0[24:5]) - temp_4));
    assign temp_7 = (((temp_3[2:1] - temp_1) != temp_1) > temp_5);
    assign temp_8 = (($unsigned(($unsigned(($signed(($unsigned(($signed(temp_4) | temp_5)) | temp_4)) | temp_4)) & temp_6[14:0])) ^ temp_2[12:3]) & temp_1);
    logic [25:0] expr_462298;
    assign expr_462298 = $signed(($signed(($signed(temp_3) * temp_6)) ^ temp_0));
    assign temp_9 = expr_462298[1:0];
    assign temp_10 = ((($unsigned((temp_6 ^ temp_7)) | temp_5) - temp_0[22:0]) ^ temp_3[2:2]);
    assign temp_11 = ($unsigned(($unsigned(($signed(($signed(($signed(temp_0) - temp_0)) != temp_6)) == (~temp_9[1:1]))) - temp_5)) <= temp_0);
    assign temp_12 = ($signed(($signed(($unsigned(($unsigned(($signed(($unsigned(temp_3[2:2]) >> input_data)) & temp_5)) & temp_2)) & temp_6)) << temp_10)) & temp_0);
    assign temp_13 = $signed(($signed(((temp_10[29:12] & temp_7) + temp_7)) ^ temp_12));
    assign temp_14 = ($unsigned(($signed((((temp_8 & temp_4) | temp_6) ^ input_data)) | temp_1)) - (~temp_5));
    assign temp_15 = (((($signed(temp_4[5:2]) >> temp_9) ^ temp_14) == temp_13[3:0]) & temp_8);
    assign temp_16 = ($signed(($unsigned(temp_13) & temp_0)) * temp_12[23:0]);
    assign temp_17 = ($signed(($unsigned(temp_3[2:0]) << temp_8)) >> temp_1[8:2]);

    assign output_data = $unsigned(($signed(((($signed(temp_6) << temp_0) + temp_10) ^ (~temp_9))) + temp_9));

endmodule