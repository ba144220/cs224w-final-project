module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;

    assign temp_0 = ($unsigned(($signed(input_data) ^ input_data)) ^ input_data);
    assign temp_1 = $signed(($unsigned(input_data) * temp_0));
    assign temp_2 = temp_1 ? ($unsigned(($unsigned((($unsigned(($unsigned(temp_0) - temp_1)) * input_data) + temp_0)) + temp_1)) + temp_0) : {3'b0, ($signed(($signed(($signed(($signed(($signed(input_data) >= temp_0)) == (~input_data))) >> temp_1)) & (~temp_0))) | temp_0)};
    assign temp_3 = temp_2;
    assign temp_4 = ($unsigned(($unsigned((($signed(($unsigned(temp_2) & (~temp_2))) * temp_0) & temp_0)) & input_data)) ^ (~temp_3));
    assign temp_5 = $unsigned(temp_0);
    assign temp_6 = ($unsigned(($unsigned(($signed(($signed(input_data[1:0]) + input_data[3:2])) & temp_1)) * input_data[2:1])) + temp_0);
    assign temp_7 = $unsigned(($signed((($unsigned((input_data | input_data)) | temp_4) * temp_0)) * temp_6));
    assign temp_8 = temp_1;
    assign temp_9 = ($signed((($unsigned(($unsigned(($signed(($unsigned((temp_1 ^ temp_4)) & temp_4)) & temp_5)) ^ temp_5)) ^ temp_4) | temp_2[30:5])) | temp_8);
    assign temp_10 = temp_4 ? ($unsigned((temp_1 ^ temp_2)) + temp_2) : $unsigned(((($unsigned(($unsigned((($signed(temp_4) - temp_9) - temp_7)) & temp_2)) * temp_6[1:1]) * temp_7) * temp_0));
    assign temp_11 = ($unsigned(($unsigned((($unsigned(((($signed(($signed((temp_5 | temp_8[18:8])) + temp_0[6:0])) ^ temp_4) - temp_8) << temp_3[7:0])) << (~temp_6)) | (~temp_10))) * temp_3)) ^ (~temp_9));

    assign output_data = ((temp_2 * temp_10[14:6]) ^ temp_2);

endmodule