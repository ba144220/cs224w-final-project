module top (
    input [3:0] input_data,
    output [36:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;
    logic [0:0] temp_13;
    logic [28:0] temp_14;
    logic [17:0] temp_15;
    logic [14:0] temp_16;
    logic [6:0] temp_17;

    assign temp_0 = 5'd13;
    assign temp_1 = ($unsigned((((temp_0 & input_data) ^ temp_0) & temp_0)) | temp_0);
    assign temp_2 = input_data;
    assign temp_3 = (($signed(temp_1) - input_data) * temp_1);
    assign temp_4 = ($signed(($unsigned(((temp_3 * temp_1) + temp_2[7:2])) - (~input_data))) + (~temp_2[7:5]));
    assign temp_5 = (($unsigned((($unsigned((temp_3 * temp_1)) | temp_0) | temp_4)) & (~temp_0)) * temp_1);
    assign temp_6 = ($signed(($signed(input_data) | temp_5[30:7])) & temp_3);
    assign temp_7 = (temp_1 ^ temp_3);
    assign temp_8 = $signed(($unsigned(($signed(($unsigned(($signed(($signed(temp_3) | input_data)) ^ input_data)) - input_data)) * temp_4)) * temp_0[4:1]));
    assign temp_9 = ((($signed((($unsigned(($signed(temp_8) * temp_5)) * temp_5) & temp_3)) & temp_4) + input_data) * temp_2);
    assign temp_10 = (($signed(($unsigned((temp_6 + temp_0)) - temp_5)) * temp_8) ^ temp_5);
    logic [31:0] expr_725303;
    assign expr_725303 = ((temp_10 ^ input_data) & temp_5);
    assign temp_11 = expr_725303[24:0];
    assign temp_12 = ($unsigned(input_data) - temp_3);
    assign temp_13 = $unsigned(($signed(($signed(temp_6) ^ input_data[1:1])) * temp_12));
    assign temp_14 = temp_2;
    logic [29:0] expr_629857;
    assign expr_629857 = ($signed(($unsigned(($unsigned(temp_8) + temp_1)) - input_data)) & temp_14);
    assign temp_15 = expr_629857[17:0];
    assign temp_16 = {10'b0, temp_0};
    assign temp_17 = (temp_6 * temp_14);

    assign output_data = ((($unsigned((temp_3[31:19] ^ temp_0)) - temp_2) | temp_10[1:0]) | (~temp_12));

endmodule