module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;
    logic [17:0] temp_12;
    logic [2:0] temp_13;
    logic [1:0] temp_14;
    logic [23:0] temp_15;
    logic [29:0] temp_16;

    assign temp_0 = (((((($signed(input_data) - input_data) | input_data) & input_data) & input_data) | input_data) * input_data);
    assign temp_1 = ((($unsigned((((($unsigned(input_data) & temp_0) + input_data) ^ temp_0) | temp_0)) ^ input_data) + temp_0[5:2]) + (~temp_0));
    assign temp_2 = $signed(($unsigned((((temp_0 * (~temp_0)) * temp_1) | temp_1)) | temp_0));
    assign temp_3 = temp_0 ? ($signed(($unsigned(($signed(($unsigned(($signed(temp_0) - temp_2[10:1])) | input_data)) ^ input_data)) | temp_0)) * temp_1) : (($signed(($signed(($unsigned(($signed(($unsigned(($unsigned(temp_2[10:1]) * temp_2)) & temp_1[23:4])) & (~input_data))) ^ temp_1[23:12])) ^ input_data)) | temp_2[10:10]) - input_data);
    assign temp_4 = $signed((($unsigned(($unsigned((((input_data + temp_3) - temp_1) - temp_0)) + temp_3)) | temp_0) ^ temp_0));
    assign temp_5 = $signed((((($signed(($signed(($signed(($unsigned((($unsigned(input_data) * (~input_data)) ^ temp_2[10:4])) * temp_3)) * temp_4)) & temp_1[16:0])) + temp_3) ^ temp_1) * temp_2) ^ temp_4));
    assign temp_6 = $unsigned((($signed(((temp_3 ^ temp_3) * input_data)) - input_data) | input_data));
    assign temp_7 = ($signed(($signed(($signed((($signed(input_data) | temp_5) & temp_1)) - temp_5)) & temp_3[19:11])) - temp_1);
    assign temp_8 = ($unsigned(($signed(($signed(($unsigned(($unsigned(($unsigned(($signed((($signed(input_data) - temp_1) & temp_7)) | temp_7)) + input_data)) - temp_4)) + temp_1)) + temp_0)) | temp_3)) - input_data);
    assign temp_9 = {4'b0, (($signed(temp_3) * temp_6) * temp_7)};
    assign temp_10 = $unsigned(($unsigned(($unsigned((temp_2 ^ temp_8[25:0])) - temp_0)) + input_data));
    assign temp_11 = ($unsigned(temp_7) ^ temp_4[16:14]);
    assign temp_12 = ($unsigned((temp_7 | temp_3)) * temp_2);
    assign temp_13 = $signed((($unsigned(($signed(temp_12) * temp_8)) ^ temp_9) ^ temp_4));
    assign temp_14 = $signed(($signed(($signed(($unsigned(temp_9) - temp_8)) & temp_7)) | temp_1));
    assign temp_15 = $signed(($signed(($unsigned(($unsigned(($unsigned(($unsigned(($signed(($unsigned(temp_3[19:2]) - temp_3)) + temp_8)) ^ temp_0)) + temp_5)) | temp_2[6:0])) | temp_13)) - temp_2[10:6]));
    assign temp_16 = ($signed(($signed(((($unsigned(($signed(temp_2) + temp_12)) | temp_13[2:2]) | temp_14) & temp_4[16:9])) ^ temp_8)) * temp_1);

    assign output_data = $signed((($unsigned(($signed(($signed(($signed(($signed(($signed(((temp_14 | temp_14) * temp_11)) ^ temp_12)) & temp_14)) * temp_5)) ^ temp_5)) * temp_10)) * temp_10) + temp_16));

endmodule