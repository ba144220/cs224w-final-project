module top (
    input [14:0] input_data,
    output [36:0] output_data
);

    logic [5:0] temp_0;
    logic [31:0] temp_1;
    logic [16:0] temp_2;
    logic [2:0] temp_3;
    logic [0:0] temp_4;
    logic [9:0] temp_5;
    logic [30:0] temp_6;

    assign temp_0 = ($signed(((((input_data[8:3] ^ (~input_data[13:8])) | input_data[9:4]) + input_data[10:5]) & input_data[12:7])) ^ input_data[9:4]);
    assign temp_1 = $unsigned(($unsigned(input_data) ^ temp_0));
    assign temp_2 = (((input_data - 17'd80248) * temp_1[14:0]) + input_data);
    assign temp_3 = temp_1;
    assign temp_4 = (temp_2 ^ input_data[6:6]);
    assign temp_5 = (((temp_3 | temp_4) - input_data[9:0]) - temp_4);
    assign temp_6 = ((temp_4 + (~temp_1)) ^ temp_0[4:0]);

    assign output_data = temp_2;

endmodule