module top (
    input [2:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;

    assign temp_0 = (((25'd27357858 & input_data) + input_data) + (~input_data));
    assign temp_1 = $signed((temp_0 & input_data));
    assign temp_2 = $signed(((input_data * temp_1) ^ input_data));
    assign temp_3 = (((temp_2[12:3] * temp_1) & input_data) + temp_2);
    logic [24:0] expr_876272;
    assign expr_876272 = temp_0;
    assign temp_4 = expr_876272[5:0];
    assign temp_5 = $unsigned(input_data);
    assign temp_6 = $unsigned(((($signed((input_data | (~input_data))) & temp_2) + input_data) | temp_5));
    assign temp_7 = $signed((((((temp_0 & temp_2) ^ input_data) + temp_2) & temp_6) ^ temp_2));
    assign temp_8 = $signed(($unsigned(((input_data | temp_6) & temp_3)) ^ temp_6));
    logic [10:0] expr_53348;
    assign expr_53348 = ((((input_data[2:1] + input_data[1:0]) + input_data[2:1]) * (~temp_1)) & temp_1);
    assign temp_9 = expr_53348[1:0];
    assign temp_10 = ((((($signed(temp_4) & temp_1) - temp_7[8:0]) & input_data) & input_data) & input_data);
    assign temp_11 = (temp_7 & (~temp_5));
    assign temp_12 = temp_7 ? ($unsigned((($signed(temp_5[8:6]) * temp_5) * input_data)) + temp_11) : (temp_7 * temp_4);
    logic [33:0] expr_714644;
    assign expr_714644 = $unsigned((($signed((($unsigned(temp_10) << (~temp_8)) | temp_10)) + (~temp_11)) * temp_10[29:7]));
    assign temp_13 = expr_714644[24:0];
    assign temp_14 = ((((temp_13 & temp_1) * temp_6) + temp_12) ^ temp_4);

    assign output_data = (temp_13 - temp_11);

endmodule