module top (
    input [5:0] input_data,
    output [5:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;

    assign temp_0 = ($unsigned(($unsigned((25'd27357858 & input_data)) + (~input_data))) + input_data);
    assign temp_1 = $signed(input_data);
    assign temp_2 = $signed(($signed(($unsigned((($unsigned(temp_1) - temp_1[8:4]) - temp_1)) ^ (~temp_0))) + temp_1));
    assign temp_3 = temp_2;
    logic [24:0] expr_876272;
    assign expr_876272 = temp_0;
    assign temp_4 = expr_876272[5:0];
    assign temp_5 = $unsigned(input_data);
    assign temp_6 = $signed(($signed(($unsigned(($signed((temp_3 & temp_5)) & temp_3)) ^ temp_0)) | temp_5));
    assign temp_7 = $signed(((temp_2[7:0] ^ temp_5) * temp_0));
    assign temp_8 = (($signed(((temp_5 | temp_1[8:5]) | temp_4)) ^ temp_5) | temp_3);
    assign temp_9 = temp_4;
    assign temp_10 = 30'd180291333;
    assign temp_11 = $unsigned(($signed((temp_0 * temp_5[2:0])) & temp_4[5:1]));
    assign temp_12 = $unsigned((($unsigned(((temp_10 ^ temp_1) - (~temp_3))) & temp_9) * temp_11));
    logic [27:0] expr_193623;
    assign expr_193623 = (($signed(temp_8) | (~temp_2)) * (~temp_4));
    assign temp_13 = expr_193623[24:0];
    assign temp_14 = (temp_9[1:1] | temp_5);

    assign output_data = $signed(($signed((temp_12 ^ temp_10[5:0])) ^ temp_5[4:0]));

endmodule