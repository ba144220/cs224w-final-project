module top (
    input [4:0] input_data,
    output [36:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;

    assign temp_0 = ($signed(input_data) ^ input_data);
    assign temp_1 = input_data[3:3] ? input_data : {5'b0, ($signed(($signed(($signed(($unsigned(($signed((($unsigned(temp_0) * temp_0) ^ temp_0)) | input_data)) ^ input_data)) | input_data)) | temp_0)) | temp_0)};
    assign temp_2 = ($unsigned((($signed(($unsigned((($unsigned(((temp_1 * temp_0) + temp_1[16:8])) - input_data) + temp_1)) + temp_1)) * temp_0) ^ temp_0)) & temp_0);
    assign temp_3 = ($signed((($signed(($unsigned(($unsigned((($unsigned((temp_1 ^ temp_0)) * temp_1) - input_data)) ^ temp_0)) - temp_2)) * temp_0) * temp_1)) & temp_2);
    assign temp_4 = ((($unsigned((temp_3 + temp_3)) * temp_3) * temp_0) + temp_0);
    assign temp_5 = ($signed(temp_0) | temp_2);
    assign temp_6 = ($unsigned(($unsigned(($signed(($unsigned((temp_2 + temp_4)) * temp_4)) & temp_4)) * temp_4)) | temp_1);

    assign output_data = ($unsigned((((($signed(temp_1) * temp_0) * temp_2) - temp_1) | temp_6)) - temp_1);

endmodule