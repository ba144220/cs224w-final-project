module top (
    input [5:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;

    assign temp_0 = (($unsigned(($unsigned(($unsigned(input_data) + input_data)) ^ (~input_data))) + input_data) | (~input_data));
    assign temp_1 = $signed(($signed(($signed((temp_0 - input_data)) & input_data)) | input_data));
    logic [27:0] expr_405099;
    assign expr_405099 = $signed((($signed(($signed(temp_0) * temp_1)) & (~temp_0)) | temp_0));
    assign temp_2 = expr_405099[12:0];
    assign temp_3 = $unsigned(3'd3);
    assign temp_4 = (($signed((($unsigned(temp_0) & input_data) - input_data)) & (~input_data)) ^ temp_0);
    assign temp_5 = (((($signed(temp_4[5:5]) * input_data) ^ temp_2) * temp_0) * temp_3);
    assign temp_6 = $unsigned(($unsigned(($signed(input_data) * temp_3)) * input_data));
    assign temp_7 = $signed(($signed(temp_1) + temp_5));
    assign temp_8 = temp_4 ? ($unsigned(((($signed(temp_0) - temp_5) - temp_5[8:2]) & (~temp_4))) | (~temp_4)) : $unsigned(($signed(input_data) + temp_1));
    assign temp_9 = ($signed(($signed(($unsigned((temp_6 * temp_7)) * temp_7)) | temp_3)) * (~temp_0));
    assign temp_10 = temp_7 ? ($unsigned(($unsigned(($signed(temp_5[8:6]) * temp_5)) * (~input_data))) - input_data) : ($unsigned(temp_7) * temp_4);
    assign temp_11 = ($unsigned(($unsigned(($unsigned(((temp_5 | (~temp_9)) ^ temp_3)) + temp_7)) ^ temp_4[5:2])) + temp_10);
    assign temp_12 = (temp_10 < temp_4);

    assign output_data = $unsigned(temp_4);

endmodule