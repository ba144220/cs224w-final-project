module top (
    input [5:0] input_data,
    output [18:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;

    assign temp_0 = ($signed(input_data) - input_data);
    assign temp_1 = (((((input_data * temp_0) * temp_0) * input_data) - input_data) | (~temp_0));
    assign temp_2 = ($signed((temp_0 | input_data)) + temp_0);
    assign temp_3 = ($unsigned(temp_2) ^ temp_2);
    assign temp_4 = $signed((($unsigned(temp_2[20:0]) * temp_2) + temp_0));
    assign temp_5 = (($signed(($unsigned(($unsigned(temp_0) - temp_1)) + temp_2)) + temp_1) - temp_4);
    assign temp_6 = ((temp_5 & temp_3[4:4]) ^ temp_5);
    assign temp_7 = ($unsigned(($signed((($unsigned(temp_0) - input_data) * temp_0)) * (~temp_6))) + temp_6);
    assign temp_8 = (temp_7 + (~temp_0[8:1]));
    assign temp_9 = $signed((($signed(temp_4) + temp_0) | temp_8));
    assign temp_10 = ((((($unsigned(temp_4) << temp_2) | temp_1) << temp_5[30:19]) & temp_0) + temp_1[4:0]);
    assign temp_11 = temp_3;
    assign temp_12 = ((((temp_10 & (~temp_9)) | temp_6) | temp_8) - temp_11);

    logic [31:0] expr_502781;
    assign expr_502781 = $signed((temp_3 * temp_10));
    assign output_data = expr_502781[18:0];

endmodule