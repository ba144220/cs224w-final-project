module top (
    input [2:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;

    assign temp_0 = (input_data + input_data);
    assign temp_1 = ((temp_0[24:8] ^ (~temp_0[24:3])) ^ temp_0);
    assign temp_2 = temp_1;
    assign temp_3 = input_data;
    assign temp_4 = (temp_2 * temp_0);
    assign temp_5 = ($unsigned(temp_1) << temp_4);
    assign temp_6 = ((temp_1[3:0] ^ temp_4) >> temp_4[5:0]);
    assign temp_7 = temp_0;
    assign temp_8 = temp_5[8:1];

    assign output_data = ((temp_5 ^ temp_8) & (~temp_8[25:20]));

endmodule