module top (
    input [3:0] input_data,
    output [18:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;
    logic [14:0] temp_13;
    logic [9:0] temp_14;
    logic [24:0] temp_15;
    logic [0:0] temp_16;
    logic [4:0] temp_17;

    assign temp_0 = input_data;
    logic [27:0] expr_753339;
    assign expr_753339 = $unsigned(((((((temp_0 - temp_0) | input_data) ^ 24'd5472715) | input_data) * temp_0) + temp_0[7:0]));
    assign temp_1 = expr_753339[23:0];
    assign temp_2 = ($signed((((($signed(((($unsigned(temp_0) | temp_0) * temp_0) ^ input_data)) | temp_0) & input_data) + input_data) ^ temp_1[2:0])) * temp_1);
    assign temp_3 = ($unsigned(temp_2) | temp_0);
    assign temp_4 = ((temp_3 + temp_1) * input_data[2:2]);
    assign temp_5 = $unsigned((($signed((((($signed(temp_3[4:4]) | input_data) ^ temp_2) * temp_1[23:0]) & temp_0)) + temp_3) | temp_0));
    logic [30:0] expr_338811;
    assign expr_338811 = temp_2;
    assign temp_6 = expr_338811[16:0];
    assign temp_7 = {6'b0, temp_0};
    assign temp_8 = (((((temp_6 - input_data) & input_data) | temp_0) ^ temp_6) + input_data);
    logic [34:0] expr_785346;
    assign expr_785346 = ($unsigned(($signed(((input_data ^ (~temp_5)) - temp_6[3:0])) & temp_0)) ^ input_data);
    assign temp_9 = expr_785346[30:0];
    assign temp_10 = temp_8 ? (temp_9 * temp_6) : ($unsigned((temp_8 & -31'd803325106)) & temp_2);
    assign temp_11 = (((((($signed(input_data) + temp_6) & input_data) ^ temp_7) + temp_3) - input_data) | temp_0);
    assign temp_12 = temp_4 ? $unsigned((($signed(((($signed(temp_7) != input_data) - temp_8) ^ temp_4)) - temp_5) != temp_11)) : ($signed(input_data) | temp_2);
    assign temp_13 = (($unsigned((((temp_2[17:0] * temp_12) + temp_1) ^ temp_11)) ^ temp_9) - temp_5);
    assign temp_14 = (($unsigned(($unsigned((temp_4 + temp_11)) - temp_7)) & temp_4) + temp_9);
    assign temp_15 = ((temp_0 * input_data) - temp_1);
    assign temp_16 = ($unsigned(temp_9[15:0]) ^ temp_5);
    assign temp_17 = ($signed(($signed((temp_6[16:13] | temp_0)) + temp_10)) + temp_7);

    assign output_data = (($signed(($unsigned((temp_14 & temp_7)) * temp_2)) ^ temp_2[17:0]) * temp_6);

endmodule