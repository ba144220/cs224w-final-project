module top (
    input [6:0] input_data,
    output [22:0] output_data
);

    logic [1:0] temp_0;
    logic [29:0] temp_1;
    logic [15:0] temp_2;
    logic [3:0] temp_3;
    logic [10:0] temp_4;
    logic [7:0] temp_5;
    logic [23:0] temp_6;
    logic [30:0] temp_7;
    logic [15:0] temp_8;
    logic [24:0] temp_9;
    logic [6:0] temp_10;

    assign temp_0 = $unsigned(input_data[4:3]);
    assign temp_1 = temp_0 ? input_data : $unsigned((temp_0 - input_data));
    assign temp_2 = ((temp_0[1:0] ^ temp_1[26:0]) + temp_0);
    assign temp_3 = ((input_data[5:2] + temp_0) | input_data[5:2]);
    logic [30:0] expr_455664;
    assign expr_455664 = (($unsigned(temp_3[3:0]) | (~temp_2)) & temp_1);
    assign temp_4 = expr_455664[10:0];
    assign temp_5 = temp_4;
    assign temp_6 = ((($signed(input_data) ^ input_data) | temp_2) ^ temp_3);
    assign temp_7 = (((temp_3 ^ temp_2) - temp_5) - temp_2);
    assign temp_8 = (((temp_4[10:3] | (~temp_2)) & input_data) & (~temp_0));
    assign temp_9 = $unsigned(((temp_1 + temp_4[9:0]) * temp_2));
    assign temp_10 = (temp_0 | temp_5);

    logic [23:0] expr_513926;
    assign expr_513926 = (((temp_2 * temp_7[30:10]) & (~temp_0[1:0])) - temp_6[18:0]);
    assign output_data = expr_513926[22:0];

endmodule