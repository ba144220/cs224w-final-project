module top (
    input [5:0] input_data,
    output [37:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;

    assign temp_0 = ($unsigned(($unsigned(($signed(input_data) & input_data)) & (~input_data))) + input_data);
    assign temp_1 = ($unsigned(($signed(((($unsigned(($unsigned(input_data) + temp_0)) | input_data) + input_data) | input_data)) * (~temp_0))) - (~temp_0));
    assign temp_2 = ($unsigned(($signed(($unsigned(($signed(temp_0[1:0]) - input_data)) * temp_0)) | temp_0)) - (~input_data));
    assign temp_3 = temp_2[21:0] ? $signed((($signed(($signed(($signed(($signed(temp_2) | temp_2[12:0])) * temp_0)) + input_data[4:0])) - temp_2) - temp_0[4:0])) : ($signed(($signed(($unsigned(temp_1) + temp_1)) ^ temp_1[23:14])) | input_data[4:0]);
    assign temp_4 = $unsigned(($unsigned(($unsigned(($signed(1'd0) ^ temp_1)) - temp_1)) * temp_3[4:2]));
    assign temp_5 = temp_2;
    assign temp_6 = temp_0 ? temp_5[17:0] : $signed((temp_2 & temp_4));

    assign output_data = temp_2;

endmodule