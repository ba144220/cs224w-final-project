module top (
    input [5:0] input_data,
    output [9:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;

    assign temp_0 = (((($unsigned(($signed(($unsigned(($unsigned((input_data | (~input_data))) | 9'd275)) ^ input_data)) - input_data)) ^ input_data) | input_data) + input_data) | input_data);
    assign temp_1 = (input_data & (~24'd13931709));
    assign temp_2 = ($unsigned(($signed(($unsigned(($unsigned(($signed(temp_0) + temp_0)) * temp_0)) | input_data)) * temp_1)) + temp_0[6:0]);
    assign temp_3 = temp_2;
    assign temp_4 = ($signed((($unsigned(($signed(($unsigned(input_data[0:0]) | input_data[4:4])) - input_data[0:0])) - temp_1[21:0]) + temp_1)) * input_data[4:4]);
    assign temp_5 = ($unsigned(((($signed(((temp_3[1:0] & input_data) ^ temp_3)) * (~input_data)) ^ (~temp_1)) ^ temp_4)) | temp_1);
    assign temp_6 = $unsigned(($signed(($unsigned(input_data) & temp_3[3:0])) + temp_0));
    assign temp_7 = (($signed(temp_4) * temp_1) * temp_5);
    assign temp_8 = ($signed((($unsigned((($signed(temp_3) | temp_6) | temp_4)) | (~temp_1)) - temp_6[3:0])) & temp_0);
    assign temp_9 = ($unsigned(temp_3[1:0]) <= temp_5);

    assign output_data = ($unsigned(($unsigned(((temp_5 & temp_8) & temp_9)) ^ temp_6)) | (~temp_7));

endmodule