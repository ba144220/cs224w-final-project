module top (
    input [3:0] input_data,
    output [9:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;
    logic [26:0] temp_10;
    logic [4:0] temp_11;
    logic [15:0] temp_12;
    logic [5:0] temp_13;
    logic [27:0] temp_14;
    logic [3:0] temp_15;
    logic [7:0] temp_16;
    logic [14:0] temp_17;

    assign temp_0 = $signed(($unsigned(($unsigned(($unsigned(($signed(input_data) + (~input_data))) * input_data)) + input_data)) | input_data));
    assign temp_1 = ($signed(($signed(input_data) + temp_0)) | input_data);
    assign temp_2 = ((temp_1 & temp_1) | temp_0);
    assign temp_3 = ($unsigned(($signed(($signed(input_data) ^ temp_1)) ^ temp_1)) | (~temp_0));
    assign temp_4 = $unsigned((($unsigned(($unsigned((($signed(($signed(temp_3) + (~input_data))) - temp_2) * temp_3)) & temp_1)) + temp_2) + input_data));
    assign temp_5 = ($unsigned(($unsigned(($unsigned(($signed(input_data) ^ (~input_data))) * temp_1)) * temp_0)) + temp_2);
    assign temp_6 = {6'b0, $signed(($unsigned((($unsigned((($signed(($signed(input_data) << input_data)) >> input_data) * temp_5)) & input_data) ^ temp_3)) << (~input_data)))};
    assign temp_7 = ($signed(temp_0) | temp_6);
    assign temp_8 = temp_3;
    assign temp_9 = ($unsigned(($signed(((($signed(input_data) & temp_1) * input_data) * temp_2)) & temp_3)) * temp_5[3:0]);
    assign temp_10 = $unsigned(input_data);
    assign temp_11 = ($unsigned((($signed(($signed(($unsigned(($signed(temp_4) | (~temp_5))) + temp_4)) * input_data)) + input_data) - temp_8)) + (~temp_8));
    assign temp_12 = $unsigned(($signed(($signed(($unsigned(($signed(($unsigned(($signed(temp_3) ^ (~temp_2))) ^ input_data)) ^ input_data)) + temp_5)) * temp_5)) + temp_1));
    assign temp_13 = ($unsigned(($signed(($unsigned(((temp_11 ^ temp_2[4:0]) - input_data)) ^ temp_11)) & temp_8)) & temp_11);
    assign temp_14 = $signed(($unsigned(temp_7) & (~input_data)));
    assign temp_15 = $unsigned((($signed(($unsigned((temp_10 & temp_8)) | temp_1)) & input_data) * input_data));
    assign temp_16 = $signed(temp_4);
    assign temp_17 = ($unsigned(($signed(($signed(temp_9) & (~temp_2))) ^ temp_4)) & (~temp_12));

    assign output_data = $signed((($signed(($unsigned(($signed((temp_17 * temp_9)) ^ temp_7)) - temp_16)) & (~temp_13)) - temp_11));

endmodule