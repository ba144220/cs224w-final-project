module top (
    input [2:0] input_data,
    output [9:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;

    assign temp_0 = ($unsigned(input_data) * input_data);
    assign temp_1 = (temp_0 | input_data);
    assign temp_2 = $unsigned(((temp_1 + temp_1) ^ temp_1));
    assign temp_3 = ($unsigned(temp_2) ^ input_data);
    assign temp_4 = temp_3;
    assign temp_5 = (temp_1[25:2] & temp_2);
    assign temp_6 = $signed(($signed((temp_0 * input_data[2:1])) - temp_1));
    assign temp_7 = (temp_6 * temp_4);
    assign temp_8 = input_data;
    assign temp_9 = ($unsigned(temp_4) & temp_4);
    assign temp_10 = {13'b0, $unsigned(temp_6)};
    assign temp_11 = $unsigned(temp_3);
    assign temp_12 = $unsigned((temp_11 * temp_2[3:0]));
    assign temp_13 = (($unsigned(temp_6) & temp_1) ^ temp_1);

    assign output_data = ($signed(temp_2) * temp_8[18:6]);

endmodule