module top (
    input [2:0] input_data,
    output [39:0] output_data
);

    logic [23:0] temp_0;
    logic [17:0] temp_1;
    logic [8:0] temp_2;
    logic [11:0] temp_3;
    logic [0:0] temp_4;
    logic [21:0] temp_5;
    logic [29:0] temp_6;
    logic [5:0] temp_7;
    logic [21:0] temp_8;
    logic [2:0] temp_9;
    logic [24:0] temp_10;
    logic [10:0] temp_11;
    logic [28:0] temp_12;
    logic [27:0] temp_13;
    logic [10:0] temp_14;
    logic [10:0] temp_15;
    logic [15:0] temp_16;
    logic [3:0] temp_17;
    logic [7:0] temp_18;

    assign temp_0 = ((input_data * input_data) + input_data);
    assign temp_1 = temp_0 ? temp_0[19:0] : ($unsigned(temp_0) <= input_data);
    assign temp_2 = input_data;
    assign temp_3 = input_data[0:0] ? temp_2 : temp_1;
    assign temp_4 = temp_2;
    assign temp_5 = temp_4 ? {6'b0, (($unsigned(temp_1[13:0]) | temp_4) + input_data)} : temp_0;
    assign temp_6 = temp_3;
    assign temp_7 = temp_4;
    assign temp_8 = ((input_data - temp_6[18:0]) | temp_0);
    logic [25:0] expr_35767;
    assign expr_35767 = ($signed(($unsigned(temp_3) ^ temp_0)) & temp_7[5:5]);
    assign temp_9 = expr_35767[2:0];
    assign temp_10 = temp_8[21:3];
    assign temp_11 = input_data[1:1] ? (temp_3 & temp_0[21:0]) : ($signed(($unsigned(temp_0) - temp_4)) * temp_5);
    assign temp_12 = (input_data + temp_3);
    assign temp_13 = temp_7 ? (temp_1 - temp_5) : ((temp_5[18:0] & temp_11) ^ temp_8);
    assign temp_14 = ($unsigned((temp_6 - temp_5)) - (~temp_12));
    assign temp_15 = temp_10;
    assign temp_16 = temp_5;
    logic [31:0] expr_371861;
    assign expr_371861 = ((temp_6 + temp_1) & temp_13);
    assign temp_17 = expr_371861[3:0];
    assign temp_18 = temp_16[11:0];

    assign output_data = temp_18;

endmodule