module top (
    input [3:0] input_data,
    output [37:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;
    logic [14:0] temp_13;

    assign temp_0 = ((((input_data | 9'd275) & input_data) & input_data) - input_data);
    assign temp_1 = {12'b0, $unsigned((((temp_0 + input_data) | input_data) * temp_0))};
    assign temp_2 = (((temp_0 | input_data) + temp_0) ^ temp_1);
    assign temp_3 = ((((input_data & temp_2) | temp_1) - temp_2) * 5'd1);
    assign temp_4 = ((input_data[3:3] + 1'd0) * temp_1);
    assign temp_5 = (temp_4 + temp_1);
    assign temp_6 = ((((temp_2 * temp_3) | input_data) ^ temp_2) * temp_1);
    assign temp_7 = temp_1;
    assign temp_8 = ((temp_0 | 13'd4485) + temp_6);
    assign temp_9 = {22'b0, temp_0};
    assign temp_10 = ((temp_6 - input_data) & temp_9);
    logic [33:0] expr_333856;
    assign expr_333856 = (((temp_5 & temp_3) & temp_0) * temp_1);
    assign temp_11 = expr_333856[25:0];
    assign temp_12 = temp_3[4:1];
    assign temp_13 = temp_1;

    assign output_data = $unsigned(temp_8[12:12]);

endmodule