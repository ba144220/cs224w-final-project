module top (
    input [2:0] input_data,
    output [36:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;

    assign temp_0 = {2'b0, input_data};
    assign temp_1 = input_data[1:1] ? ((temp_0 | temp_0) & input_data) : (input_data * temp_0);
    assign temp_2 = input_data;
    assign temp_3 = ((input_data ^ input_data) - input_data);
    assign temp_4 = {10'b0, ((temp_1 & input_data) | temp_2[7:5])};
    assign temp_5 = temp_4;
    assign temp_6 = input_data;
    assign temp_7 = input_data;
    assign temp_8 = temp_4;
    assign temp_9 = temp_2;
    logic [17:0] expr_921402;
    assign expr_921402 = ((temp_0 * temp_6[10:0]) + temp_1);
    assign temp_10 = expr_921402[1:0];
    assign temp_11 = ((temp_2 ^ temp_0) & temp_7);

    assign output_data = temp_9;

endmodule