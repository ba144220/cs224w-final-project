module top (
    input [4:0] input_data,
    output [16:0] output_data
);

    logic [22:0] temp_0;
    logic [1:0] temp_1;
    logic [29:0] temp_2;
    logic [15:0] temp_3;
    logic [3:0] temp_4;
    logic [10:0] temp_5;
    logic [7:0] temp_6;
    logic [23:0] temp_7;
    logic [30:0] temp_8;
    logic [15:0] temp_9;
    logic [24:0] temp_10;

    assign temp_0 = (((($unsigned(input_data) & input_data) + input_data) - input_data) ^ input_data);
    assign temp_1 = $unsigned(($unsigned((temp_0 + temp_0)) - temp_0));
    assign temp_2 = temp_0;
    assign temp_3 = (($unsigned(((temp_1[1:1] - temp_2) + temp_1)) * input_data) + temp_2);
    assign temp_4 = ((temp_1 + temp_2) | input_data[4:1]);
    assign temp_5 = (temp_1 * temp_3);
    assign temp_6 = temp_2;
    assign temp_7 = ($unsigned((temp_4 * temp_6)) * temp_6);
    assign temp_8 = (temp_4 ^ temp_6);
    assign temp_9 = ((((temp_0 - temp_2) & temp_6[7:2]) + temp_4) + temp_4);
    assign temp_10 = ((((temp_9 - temp_9) * temp_9) & temp_3) - (~temp_4));

    assign output_data = (temp_9 + temp_2[29:18]);

endmodule