module top (
    input [3:0] input_data,
    output [37:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;

    assign temp_0 = (((input_data & (~input_data)) | (~input_data)) | 9'd275);
    assign temp_1 = ((((((input_data + temp_0) * temp_0) * input_data) - input_data) | (~temp_0)) + (~temp_0));
    assign temp_2 = $unsigned((((((temp_0 + temp_0) ^ temp_1) & input_data) | temp_0) * temp_1));
    assign temp_3 = $unsigned(((((($signed(temp_2) * temp_1) | temp_1) - temp_0) ^ temp_0) - temp_2));
    assign temp_4 = ((1'd0 & temp_2) + input_data[0:0]);
    assign temp_5 = (((temp_4 & (~temp_4)) != (~temp_1)) != temp_4);
    assign temp_6 = ($unsigned(($signed(((temp_0 | temp_0) + temp_4)) | (~temp_0))) + temp_3);

    assign output_data = ($signed(($signed(($unsigned(($signed(temp_2[30:1]) ^ temp_5[30:6])) | temp_3[4:4])) * temp_3)) | temp_0);

endmodule