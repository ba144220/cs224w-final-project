module top (
    input [9:0] input_data,
    output [39:0] output_data
);

    logic [23:0] temp_0;
    logic [17:0] temp_1;
    logic [8:0] temp_2;
    logic [11:0] temp_3;
    logic [0:0] temp_4;
    logic [21:0] temp_5;
    logic [29:0] temp_6;
    logic [5:0] temp_7;
    logic [21:0] temp_8;
    logic [2:0] temp_9;
    logic [24:0] temp_10;
    logic [10:0] temp_11;
    logic [28:0] temp_12;
    logic [27:0] temp_13;
    logic [10:0] temp_14;

    assign temp_0 = input_data;
    assign temp_1 = $signed((temp_0 - temp_0));
    assign temp_2 = temp_0[23:19] ? (((temp_0 | temp_1) + input_data[8:0]) | input_data[8:0]) : temp_0;
    assign temp_3 = (((temp_2 - temp_1) + temp_2) ^ temp_2);
    assign temp_4 = ((temp_1 + temp_0[15:0]) | temp_2);
    logic [28:0] expr_632205;
    assign expr_632205 = ((((((input_data ^ (~temp_4)) | temp_0) & temp_4) * temp_0) | (~temp_0)) - input_data);
    assign temp_5 = expr_632205[21:0];
    assign temp_6 = temp_3 ? (((((((temp_4 - temp_0) >> temp_3[2:0]) + temp_3) - input_data) & temp_0) + (~temp_4)) & temp_2[8:2]) : (((((((temp_0 + input_data) * 30'd530821750) | temp_3) | temp_3) | temp_1) * input_data) * temp_5);
    assign temp_7 = $signed(temp_0);
    assign temp_8 = ((((((input_data | temp_5) | temp_2[8:1]) ^ temp_1) - temp_2) * temp_2) * temp_2);
    assign temp_9 = $unsigned((((((temp_6 & temp_2) >> input_data[2:0]) & input_data[2:0]) & (~temp_5)) << temp_3));
    assign temp_10 = $unsigned(((((((input_data + input_data) ^ temp_1) * temp_3) + temp_0) + temp_6) - temp_0));
    assign temp_11 = (temp_2 | temp_6);
    assign temp_12 = input_data[7:7] ? $signed(((((temp_11 * temp_10) & temp_11) & temp_4) & temp_0)) : (input_data | temp_4);
    assign temp_13 = (((((temp_0 & temp_1) & temp_8) & temp_9) | temp_12) ^ temp_8);
    assign temp_14 = $signed((((((temp_11 | temp_12) - temp_13) ^ temp_9) + temp_4) * temp_1));

    assign output_data = (((temp_6 & temp_3) ^ temp_2) + temp_9);

endmodule