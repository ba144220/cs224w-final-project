module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;

    assign temp_0 = $signed(input_data);
    assign temp_1 = $signed((input_data - temp_0));
    assign temp_2 = $signed(((temp_1 + temp_1) * temp_0[2:0]));
    assign temp_3 = temp_0;
    assign temp_4 = (input_data ^ input_data);
    assign temp_5 = $unsigned(((temp_3 | input_data) * input_data));
    assign temp_6 = $signed(((temp_0 * input_data[3:2]) ^ input_data[1:0]));
    assign temp_7 = temp_1;
    assign temp_8 = (temp_6 != temp_7);
    assign temp_9 = (input_data * input_data);
    assign temp_10 = (($unsigned(temp_0) & (~temp_6)) * temp_6);
    assign temp_11 = $unsigned((temp_9[3:0] * temp_2[3:0]));
    assign temp_12 = ((input_data & temp_1) & temp_7[7:0]);
    logic [26:0] expr_257363;
    assign expr_257363 = (temp_7 + temp_0[6:1]);
    assign temp_13 = expr_257363[11:0];
    assign temp_14 = (input_data | temp_8);
    assign temp_15 = (temp_10 | temp_12);

    assign output_data = $unsigned(temp_5);

endmodule