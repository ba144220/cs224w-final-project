module top (
    input [2:0] input_data,
    output [18:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;
    logic [14:0] temp_13;
    logic [9:0] temp_14;
    logic [24:0] temp_15;
    logic [0:0] temp_16;
    logic [4:0] temp_17;
    logic [10:0] temp_18;

    assign temp_0 = {8'b0, ((input_data > input_data) < input_data)};
    assign temp_1 = (temp_0 | temp_0);
    assign temp_2 = temp_0;
    assign temp_3 = temp_1;
    assign temp_4 = temp_2;
    assign temp_5 = temp_1;
    assign temp_6 = (input_data | temp_4);
    assign temp_7 = ($unsigned(temp_2[14:0]) | temp_3);
    assign temp_8 = $unsigned(((13'd7476 * temp_5[6:0]) | temp_6[1:0]));
    assign temp_9 = ($unsigned(temp_1) ^ temp_7);
    assign temp_10 = temp_9;
    assign temp_11 = ($signed((temp_4 * (~temp_6[14:0]))) | input_data);
    assign temp_12 = 10'd71;
    assign temp_13 = temp_0;
    assign temp_14 = temp_0 ? (temp_12 - temp_13[4:0]) : temp_12;
    assign temp_15 = (temp_12[2:0] + temp_0);
    assign temp_16 = (($signed(input_data[0:0]) | temp_12) | temp_1);
    assign temp_17 = (temp_2 * temp_10);
    assign temp_18 = $signed(((temp_3 + temp_0) | temp_12[1:0]));

    assign output_data = ((temp_2[25:0] | temp_16) | temp_1);

endmodule