module top (
    input [4:0] input_data,
    output [18:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;
    logic [0:0] temp_13;
    logic [28:0] temp_14;
    logic [17:0] temp_15;

    assign temp_0 = $unsigned(input_data);
    assign temp_1 = (input_data & input_data);
    assign temp_2 = ((input_data != input_data) & (~temp_1));
    assign temp_3 = input_data;
    assign temp_4 = ($signed((input_data ^ input_data)) - input_data);
    assign temp_5 = ((input_data & temp_0) << temp_2[7:5]);
    assign temp_6 = temp_4;
    assign temp_7 = input_data;
    assign temp_8 = input_data;
    assign temp_9 = input_data;
    logic [26:0] expr_313111;
    assign expr_313111 = (($unsigned(temp_6) - temp_8) | temp_8);
    assign temp_10 = expr_313111[1:0];
    assign temp_11 = input_data;
    assign temp_12 = temp_3;
    assign temp_13 = (($unsigned(temp_1) << (~temp_7[11:0])) << temp_0);
    assign temp_14 = temp_13;
    assign temp_15 = temp_4;

    assign output_data = ($unsigned(temp_15) + temp_10[1:0]);

endmodule