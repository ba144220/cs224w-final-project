module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;

    assign temp_0 = ($unsigned((($signed(($unsigned((input_data + input_data)) * input_data)) | input_data) | input_data)) * input_data);
    assign temp_1 = input_data;
    assign temp_2 = ($signed(temp_1) | temp_0[6:1]);
    assign temp_3 = ($signed((($unsigned(($unsigned(temp_1) + temp_1)) - (~temp_0)) + temp_1[12:0])) >> input_data);
    assign temp_4 = ($signed(($unsigned(((($unsigned(($signed(($signed(temp_2) - temp_1)) & temp_3[9:5])) * temp_0) ^ temp_0[6:2]) - temp_3)) ^ temp_2)) ^ temp_0);
    assign temp_5 = $unsigned(($unsigned((($signed((($signed(($signed((temp_0[6:5] * temp_3)) ^ (~temp_4))) | temp_4) | (~input_data))) | temp_1) + temp_4)) ^ temp_0));
    assign temp_6 = ($unsigned(($unsigned(temp_0[6:3]) + temp_3)) * temp_1);
    assign temp_7 = (($unsigned(($unsigned(($signed(temp_4[5:5]) * input_data)) - (~temp_2))) ^ temp_1) | input_data);
    assign temp_8 = (temp_7 | temp_4);
    assign temp_9 = ($signed((($unsigned(($unsigned((temp_6 * temp_6)) | temp_5)) ^ temp_4) | (~temp_2[30:5]))) | temp_8);

    assign output_data = temp_4[3:0] ? ($unsigned(($unsigned(temp_2) | (~temp_5))) * temp_7) : ($unsigned((($unsigned(($unsigned(($unsigned(($signed(temp_6) ^ temp_0)) + temp_3[9:9])) ^ temp_6[1:1])) * temp_6[1:1]) * temp_7)) * temp_1);

endmodule