module top (
    input [4:0] input_data,
    output [18:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;

    assign temp_0 = input_data;
    assign temp_1 = temp_0 ? $signed((($unsigned((input_data | temp_0)) & input_data) + input_data)) : $unsigned(((((((($unsigned(17'd105981) & (~input_data)) - input_data) * (~input_data)) - input_data) | temp_0) ^ (~17'd53866)) * input_data));
    assign temp_2 = ((((($unsigned((($unsigned(input_data) + (~input_data)) + temp_1)) + temp_1) * (~temp_0)) + temp_0) & temp_0) ^ (~input_data));
    assign temp_3 = ((($signed(($signed(((input_data - input_data) | temp_2)) >= temp_2)) < temp_1) < 32'd3361672518) == temp_1);
    assign temp_4 = input_data;
    assign temp_5 = $unsigned(($signed(((($unsigned((input_data - temp_0)) - input_data) * temp_2) + 31'd393776021)) + temp_4));
    assign temp_6 = {4'b0, $unsigned(($unsigned(($unsigned(($signed((temp_1 + input_data)) + temp_2)) | input_data)) - temp_2))};
    assign temp_7 = ((((temp_6 + (~input_data)) + temp_0) - (~temp_6)) - input_data);
    assign temp_8 = temp_0 ? (((temp_3 & temp_4) * temp_7) + temp_2) : (temp_7 & temp_7);
    assign temp_9 = (((temp_5 & temp_4) >= (~temp_1)) | temp_0);
    assign temp_10 = (temp_1 | temp_1);
    assign temp_11 = temp_2 ? $signed((((temp_1 & (~temp_0)) | temp_4) | (~temp_10))) : (((temp_1 | temp_8) + temp_9) * temp_7);

    assign output_data = temp_6 ? ($unsigned((((temp_11 & temp_9) * temp_11) + temp_10)) | temp_11) : {17'b0, $signed(temp_10)};

endmodule