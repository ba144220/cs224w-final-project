module top (
    input [3:0] input_data,
    output [2:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;

    assign temp_0 = input_data;
    assign temp_1 = temp_0;
    assign temp_2 = $unsigned((($unsigned(((($signed(temp_0) - input_data) | temp_0) | temp_0)) == temp_1) > temp_1));
    assign temp_3 = $unsigned((((($unsigned(((($signed((($signed(temp_0[6:3]) ^ temp_1) ^ temp_2[30:20])) - temp_2) * input_data) - temp_0[2:0])) | temp_1) & (~temp_0)) & (~temp_2)) * temp_2));
    assign temp_4 = $unsigned(((((((temp_0[6:2] | temp_1) & temp_2) * input_data) * temp_0) & input_data) | temp_0));
    assign temp_5 = (((((($unsigned(($unsigned((temp_0[6:0] | temp_4)) | temp_2)) * temp_3) * temp_3) - temp_3) - temp_2) ^ temp_2[30:26]) + temp_3);
    assign temp_6 = ((($unsigned(((temp_4 & temp_3) * temp_0)) * temp_2) * temp_2) + temp_0);
    assign temp_7 = $signed((temp_1 | temp_5));
    assign temp_8 = (((((((temp_5 + temp_7) | temp_1) * temp_4) + temp_3[3:0]) | temp_4[2:0]) + temp_1[25:21]) ^ temp_2);

    assign output_data = (((((($signed(((temp_3 - temp_6) == temp_4)) + temp_4[5:2]) + temp_3[9:9]) != temp_6) > temp_5) + temp_3) > temp_5[4:2]);

endmodule