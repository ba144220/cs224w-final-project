module top (
    input [3:0] input_data,
    output [37:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;
    logic [14:0] temp_13;
    logic [9:0] temp_14;
    logic [24:0] temp_15;

    assign temp_0 = (((((input_data * input_data) & input_data) & (~input_data)) - input_data) ^ input_data);
    logic [27:0] expr_628896;
    assign expr_628896 = (($unsigned(($unsigned((24'd5472715 ^ input_data)) | temp_0[8:0])) - (~temp_0)) ^ input_data);
    assign temp_1 = expr_628896[23:0];
    assign temp_2 = (temp_0 * input_data);
    assign temp_3 = temp_1;
    assign temp_4 = ((temp_2[20:0] * temp_2) >> temp_0);
    assign temp_5 = (input_data + 31'd564447966);
    assign temp_6 = (((temp_2 - temp_5) + temp_1) * input_data);
    assign temp_7 = ((((($signed(temp_3[4:4]) | input_data) ^ temp_2) * temp_1[23:0]) & temp_0) + temp_3[1:0]);
    assign temp_8 = ((input_data * input_data) & (~temp_4));
    assign temp_9 = (temp_0 <= temp_2);
    assign temp_10 = temp_1;
    assign temp_11 = (((((temp_5 * temp_6) + temp_3) | temp_4) | temp_10) ^ temp_2);
    assign temp_12 = ((temp_10 * temp_1[19:0]) + temp_1);
    assign temp_13 = (input_data * temp_1);
    assign temp_14 = $signed(($signed((((temp_10 - temp_11) - temp_12) ^ temp_12)) | input_data));
    assign temp_15 = {9'b0, (temp_3 ^ temp_7)};

    assign output_data = $unsigned((temp_2 - temp_6));

endmodule