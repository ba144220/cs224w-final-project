module top (
    input [2:0] input_data,
    output [31:0] output_data
);

    logic [16:0] temp_0;
    logic [2:0] temp_1;
    logic [0:0] temp_2;
    logic [9:0] temp_3;
    logic [30:0] temp_4;
    logic [23:0] temp_5;
    logic [20:0] temp_6;
    logic [1:0] temp_7;
    logic [17:0] temp_8;
    logic [31:0] temp_9;
    logic [12:0] temp_10;
    logic [26:0] temp_11;

    assign temp_0 = (($signed(((input_data ^ input_data) + input_data)) + input_data) ^ input_data);
    assign temp_1 = (((($signed(temp_0) - temp_0) * temp_0[16:11]) | temp_0) << temp_0);
    assign temp_2 = $unsigned(input_data[0:0]);
    assign temp_3 = (temp_1 ^ input_data);
    assign temp_4 = (((temp_3 | temp_2) * temp_3[9:2]) & 31'd1156433848);
    assign temp_5 = (($unsigned(($signed(input_data) | temp_0[16:4])) + temp_4) ^ temp_0[16:7]);
    assign temp_6 = ($signed((((input_data + temp_2) + (~temp_1)) - temp_0)) ^ temp_0);
    assign temp_7 = temp_5;
    assign temp_8 = ($signed(($signed((($signed(temp_5) + temp_6) | temp_2)) ^ (~temp_2))) + temp_1);
    assign temp_9 = temp_2;
    assign temp_10 = temp_4;
    assign temp_11 = ($unsigned(temp_10) + temp_1);

    assign output_data = temp_0;

endmodule