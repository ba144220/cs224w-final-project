module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;

    assign temp_0 = input_data;
    assign temp_1 = ($signed(($signed(temp_0) + input_data)) * input_data);
    assign temp_2 = temp_1;
    assign temp_3 = ($unsigned(($signed(($signed(($unsigned(($unsigned(temp_2) - -10'd118)) + temp_0[6:3])) ^ temp_1[10:0])) | temp_0)) - temp_0);
    assign temp_4 = ($signed(temp_1) & temp_0);
    assign temp_5 = $signed(temp_3);
    assign temp_6 = ($signed(temp_2) & (~input_data[3:2]));
    assign temp_7 = ($signed(temp_5) - temp_5);
    assign temp_8 = ($unsigned(($signed((input_data * temp_7)) + temp_2[29:0])) << input_data);
    assign temp_9 = (($signed(($signed(temp_7) << (~temp_5[1:0]))) <= temp_3) - temp_5);
    assign temp_10 = ($signed(($unsigned(temp_8) - temp_5)) + (~temp_1));
    assign temp_11 = ($unsigned(temp_9) & temp_9);
    assign temp_12 = ($signed(($unsigned(($unsigned(($unsigned(($unsigned(temp_10) * temp_5)) * temp_5)) + temp_1)) + temp_7)) ^ temp_9);
    assign temp_13 = (((temp_7[25:6] | temp_8) - temp_7) * temp_12);
    assign temp_14 = ($unsigned((temp_9 | (~temp_3[9:1]))) | temp_10);
    assign temp_15 = (($unsigned(($unsigned((temp_2 | temp_1)) | temp_5[4:1])) * temp_1) * temp_7);
    assign temp_16 = ($signed(((($unsigned(temp_11) & temp_1) & temp_10[14:4]) ^ temp_1)) + temp_1);

    assign output_data = (($signed((($unsigned(($unsigned(temp_16[13:4]) | temp_8[18:2])) - (~temp_11)) & temp_15)) ^ (~temp_9)) & temp_8);

endmodule