module top (
    input [5:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;

    assign temp_0 = ($unsigned((input_data + input_data)) ^ input_data);
    assign temp_1 = temp_0 ? temp_0 : ((input_data - temp_0) & input_data);
    assign temp_2 = ((input_data * temp_1) & (~temp_0));
    assign temp_3 = (input_data[2:0] | temp_2[2:0]);
    logic [25:0] expr_911111;
    assign expr_911111 = ($unsigned(temp_0) ^ temp_2);
    assign temp_4 = expr_911111[5:0];
    assign temp_5 = $signed((($unsigned(temp_0[20:0]) - temp_3) ^ temp_0));
    assign temp_6 = ($unsigned((input_data | temp_5)) - temp_3);
    assign temp_7 = temp_5;
    assign temp_8 = (input_data & input_data);
    assign temp_9 = ((temp_5 | temp_1) & temp_4);
    assign temp_10 = temp_3;
    assign temp_11 = temp_9;
    assign temp_12 = ($signed((temp_10 - (~temp_5))) - (~temp_10));

    assign output_data = (temp_11 - (~temp_4));

endmodule