module top (
    input [3:0] input_data,
    output [37:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;

    assign temp_0 = (($unsigned(($signed(input_data) & input_data)) & (~input_data)) + input_data);
    assign temp_1 = ($unsigned(($unsigned(((((input_data + temp_0) * temp_0) * temp_0) * input_data)) | temp_0[8:0])) - (~temp_0));
    assign temp_2 = ($signed(((($signed(temp_0) - input_data) * temp_0) ^ input_data)) | temp_0);
    assign temp_3 = $unsigned(((((($signed((temp_2 * (~temp_1[23:2]))) * temp_1) | temp_1) - temp_0) ^ temp_0) - temp_2));
    assign temp_4 = $unsigned((($signed(($signed(($unsigned(((((((($signed((($unsigned(temp_0) - (~temp_2)) & temp_0)) | input_data[1:1]) ^ temp_2) * temp_1[23:0]) & temp_0) + temp_3[1:0]) | temp_0) - (~temp_2))) ^ temp_3[3:0])) + temp_0)) + temp_0) & (~temp_2)));
    assign temp_5 = $unsigned(temp_3[4:4]);

    assign output_data = $unsigned(((($signed(((((($signed(((($signed(temp_1) + temp_3) | temp_2) | (~temp_3))) | temp_5[5:0]) | temp_0) + temp_0) | temp_2[30:25]) - temp_0)) | temp_1) & temp_2) + temp_3));

endmodule