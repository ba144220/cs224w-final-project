module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;

    logic [7:0] expr_48572;
    assign expr_48572 = $unsigned(((((((input_data | input_data) + input_data) | input_data) << input_data) | 7'd79) << input_data));
    assign temp_0 = input_data[2:2] ? expr_48572[6:0] : $signed((((input_data ^ input_data) ^ input_data) | input_data));
    assign temp_1 = ((((input_data + temp_0) + temp_0) - temp_0) * temp_0);
    assign temp_2 = $unsigned((temp_0 - temp_1));
    assign temp_3 = $unsigned((temp_1 & temp_1[25:9]));
    assign temp_4 = temp_0 ? $unsigned((((((temp_3 | temp_1) & temp_2) * temp_1[20:0]) ^ temp_1) & temp_0)) : (temp_2 & temp_3[1:0]);

    assign output_data = $signed(temp_4);

endmodule