module top (
    input [2:0] input_data,
    output [9:0] output_data
);

    logic [23:0] temp_0;
    logic [17:0] temp_1;
    logic [8:0] temp_2;
    logic [11:0] temp_3;
    logic [0:0] temp_4;
    logic [21:0] temp_5;
    logic [29:0] temp_6;
    logic [5:0] temp_7;
    logic [21:0] temp_8;
    logic [2:0] temp_9;
    logic [24:0] temp_10;
    logic [10:0] temp_11;

    assign temp_0 = $unsigned((((((((input_data + input_data) ^ input_data) & input_data) * input_data) & 24'd16499108) ^ input_data) | input_data));
    assign temp_1 = $unsigned(((((((((temp_0 | 18'd78278) | input_data) | input_data) | temp_0) | temp_0) * 18'd13312) & input_data) ^ temp_0));
    assign temp_2 = input_data[1:1] ? $unsigned(((temp_0 * input_data) * temp_0)) : $signed((((((((((input_data * temp_0) - input_data) | input_data) * input_data) & input_data) * temp_0) & input_data) - temp_1) ^ temp_0[2:0]));
    assign temp_3 = temp_1[15:0];
    assign temp_4 = ((temp_1 - temp_0) > input_data[2:2]);
    assign temp_5 = temp_0;
    assign temp_6 = (((temp_0 & input_data) * temp_3) & temp_0);
    assign temp_7 = (((((temp_1 * 6'd49) ^ temp_5) <= temp_3) + input_data) - temp_6);
    assign temp_8 = (((((input_data | temp_4) ^ temp_1) - temp_2) * temp_2) * temp_2);
    assign temp_9 = temp_0;
    assign temp_10 = (((25'd16583682 & input_data) ^ temp_2[4:0]) ^ temp_4);
    assign temp_11 = $unsigned(((temp_8 | temp_6[13:0]) ^ temp_10));

    assign output_data = temp_10;

endmodule