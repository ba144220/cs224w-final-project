module top (
    input [2:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;

    assign temp_0 = ($unsigned(input_data) + input_data);
    assign temp_1 = input_data;
    assign temp_2 = ($signed(($unsigned(input_data) & input_data)) * input_data);
    logic [10:0] expr_695385;
    assign expr_695385 = (($signed(temp_1) | input_data) * temp_1);
    assign temp_3 = expr_695385[2:0];
    assign temp_4 = temp_0;
    assign temp_5 = $unsigned(temp_4[1:0]);
    assign temp_6 = temp_4[1:0];
    assign temp_7 = $unsigned(14'd6883);
    assign temp_8 = {11'b0, $signed(($signed(($unsigned(temp_1[4:0]) & temp_2)) | temp_7))};
    assign temp_9 = temp_8;

    assign output_data = $signed(($unsigned(($unsigned(temp_9) ^ temp_6)) ^ temp_8));

endmodule