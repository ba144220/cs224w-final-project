module top (
    input [3:0] input_data,
    output [18:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;
    logic [0:0] temp_13;
    logic [28:0] temp_14;
    logic [17:0] temp_15;

    assign temp_0 = $unsigned(input_data);
    assign temp_1 = temp_0;
    assign temp_2 = (input_data - temp_1);
    assign temp_3 = $unsigned(($unsigned((input_data | input_data)) | input_data));
    assign temp_4 = (input_data == temp_1);
    assign temp_5 = $unsigned(((temp_4[28:26] ^ temp_1) * temp_1));
    assign temp_6 = $signed((($unsigned(temp_4) <= input_data) + temp_2));
    assign temp_7 = (temp_3[31:13] * temp_1);
    assign temp_8 = temp_2;
    assign temp_9 = {5'b0, ((temp_0 * temp_6) * temp_1)};
    assign temp_10 = input_data[3:2];
    assign temp_11 = temp_6;
    assign temp_12 = $signed(((temp_4[7:0] * temp_9) & input_data));
    assign temp_13 = ((temp_4 * temp_9) + temp_6);
    assign temp_14 = $signed(($signed(temp_4) <= temp_7));
    assign temp_15 = $unsigned(temp_1);

    assign output_data = ((temp_8 - temp_10[1:1]) & temp_10);

endmodule