module top (
    input [2:0] input_data,
    output [9:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;
    logic [1:0] temp_17;

    assign temp_0 = ($unsigned((input_data + input_data)) - input_data);
    assign temp_1 = ((temp_0 * temp_0[4:0]) | input_data);
    assign temp_2 = ((input_data * temp_0) + temp_0[6:3]);
    assign temp_3 = temp_2;
    assign temp_4 = (temp_1[25:2] & temp_2);
    assign temp_5 = (temp_4 + temp_4);
    assign temp_6 = (input_data[2:1] - temp_2);
    assign temp_7 = ((temp_5 ^ temp_3[4:0]) - temp_5);
    logic [32:0] expr_918996;
    assign expr_918996 = ((temp_4 + temp_2) ^ (~temp_7));
    assign temp_8 = expr_918996[18:0];
    assign temp_9 = ($unsigned(((input_data - temp_5) & temp_0)) - temp_1);
    assign temp_10 = ((input_data + input_data) ^ temp_1);
    logic [27:0] expr_55490;
    assign expr_55490 = (($unsigned(temp_7) + temp_0) | temp_3);
    assign temp_11 = expr_55490[23:0];
    assign temp_12 = ((temp_9 & temp_7) * temp_1);
    assign temp_13 = input_data;
    assign temp_14 = temp_12 ? temp_9 : (temp_9 ^ temp_9);
    assign temp_15 = (((temp_13 | temp_2) & input_data) ^ temp_9);
    assign temp_16 = temp_1;
    assign temp_17 = ((temp_6[1:0] - temp_1) * temp_13);

    assign output_data = (((temp_15 - temp_8) - temp_12[1:0]) * temp_4[1:0]);

endmodule