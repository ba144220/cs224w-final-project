module top (
    input [3:0] input_data,
    output [37:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;

    assign temp_0 = (((((((((((input_data - input_data) + (~input_data)) * input_data) & (~input_data)) * input_data) ^ input_data) | input_data) ^ input_data) ^ input_data) | input_data) * input_data);
    assign temp_1 = ((temp_0[1:0] < input_data) | temp_0[8:4]);
    assign temp_2 = ($signed(((((input_data | temp_0) ^ input_data) | temp_1) - temp_1)) ^ temp_0[8:6]);
    assign temp_3 = $signed((((((input_data | temp_0) - temp_2) - temp_0[4:0]) - 5'd20) - input_data));
    assign temp_4 = (((((temp_0 + (~temp_3)) & input_data[2:2]) + (~input_data[0:0])) ^ (~temp_1)) ^ temp_2[30:18]);
    assign temp_5 = ($signed((($unsigned(((((($signed((($signed(($signed(($unsigned((temp_1 + (~temp_2))) ^ temp_3[3:0])) + temp_0)) + temp_0) & (~temp_2))) + temp_3) | temp_0) ^ temp_3) + temp_1) | temp_2)) | (~temp_0)) - temp_3[1:0])) & temp_0);
    assign temp_6 = ($signed(temp_5) - temp_0);
    assign temp_7 = ((((((temp_4 | temp_3) | temp_4) - temp_5) - temp_6) ^ temp_6) | temp_1);

    assign output_data = (((((($unsigned(($signed((($signed(($signed(($signed(($unsigned((temp_7 | temp_0)) ^ temp_0)) - temp_4)) + temp_4)) + temp_1) * temp_0[6:0])) - temp_7)) + temp_7) * temp_7) * temp_1) + temp_7[14:5]) - (~temp_2)) | temp_2);

endmodule