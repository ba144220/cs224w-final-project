module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;

    assign temp_0 = ($unsigned(($signed(input_data) ^ input_data)) ^ input_data);
    assign temp_1 = ($unsigned(input_data) * temp_0);
    assign temp_2 = input_data;
    assign temp_3 = ($unsigned(temp_1) | temp_2);
    assign temp_4 = ($unsigned(($unsigned(temp_0) ^ temp_2)) - temp_1);
    assign temp_5 = ($unsigned(($signed(($signed(($unsigned(($signed(temp_0) - (~temp_0))) & temp_2)) - temp_1)) & temp_3[9:5])) * temp_0);
    assign temp_6 = temp_4;
    assign temp_7 = ($unsigned(($unsigned(($signed(($signed(($unsigned(temp_5) & 26'd25670156)) * temp_0)) & temp_0)) & temp_4)) | temp_3);
    assign temp_8 = $unsigned(temp_0);
    assign temp_9 = ($unsigned(($signed(($unsigned(($unsigned(temp_6) | (~temp_5))) - temp_7)) - temp_5)) + temp_7);
    assign temp_10 = temp_7;
    logic [31:0] expr_192825;
    assign expr_192825 = ($unsigned(($signed(($unsigned((($unsigned(($unsigned(($unsigned(temp_10) | temp_9)) | temp_1)) * temp_9) + temp_9)) + temp_7)) ^ temp_9)) | temp_7);
    assign temp_11 = expr_192825[23:0];

    assign output_data = $unsigned(($signed(($unsigned((($unsigned(($signed(($signed((temp_5 + temp_2)) * temp_9)) & temp_9)) - temp_6) | temp_3[9:1])) * temp_0)) - temp_10));

endmodule