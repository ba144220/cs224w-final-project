module top (
    input [3:0] input_data,
    output [31:0] output_data
);

    logic [16:0] temp_0;
    logic [2:0] temp_1;
    logic [0:0] temp_2;
    logic [9:0] temp_3;
    logic [30:0] temp_4;
    logic [23:0] temp_5;
    logic [20:0] temp_6;
    logic [1:0] temp_7;
    logic [17:0] temp_8;
    logic [31:0] temp_9;

    assign temp_0 = ($signed(((input_data ^ input_data) + input_data)) + input_data);
    assign temp_1 = $unsigned(($unsigned(input_data[2:0]) ^ temp_0));
    assign temp_2 = (((input_data[0:0] - 1'd1) * temp_1) & temp_0);
    assign temp_3 = (((input_data & temp_0[4:0]) - temp_1) & temp_1);
    assign temp_4 = ((input_data * temp_3) | temp_0);
    assign temp_5 = temp_0;
    assign temp_6 = {19'b0, temp_1[2:1]};
    assign temp_7 = temp_6;
    assign temp_8 = (((temp_3 >> temp_4) ^ temp_0) << temp_5[3:0]);
    assign temp_9 = ((temp_3 - (~temp_1[2:2])) ^ temp_0);

    assign output_data = (temp_2 * temp_3[9:7]);

endmodule