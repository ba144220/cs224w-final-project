module top (
    input [2:0] input_data,
    output [31:0] output_data
);

    logic [16:0] temp_0;
    logic [2:0] temp_1;
    logic [0:0] temp_2;
    logic [9:0] temp_3;
    logic [30:0] temp_4;
    logic [23:0] temp_5;

    assign temp_0 = input_data;
    assign temp_1 = ($signed((((temp_0 & input_data) * temp_0) - temp_0)) + temp_0);
    assign temp_2 = temp_1;
    assign temp_3 = ((temp_1 | temp_1) & temp_1);
    assign temp_4 = temp_2 ? ((((temp_3 & temp_3) ^ temp_2) ^ temp_2) * temp_3) : {11'b0, (($unsigned(((($unsigned((($unsigned(temp_2) >> temp_1) * temp_0)) - temp_1) >> temp_0) >> (~temp_3))) | input_data) >> temp_2)};
    assign temp_5 = $unsigned((((((temp_1 - temp_0) * temp_4) != temp_4) != temp_3) + temp_4));

    assign output_data = $signed((($signed(temp_5) - temp_1) + temp_0));

endmodule