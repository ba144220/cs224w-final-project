module top (
    input [5:0] input_data,
    output [37:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;

    assign temp_0 = ((((((input_data != 9'd163) | input_data) < input_data) > (~input_data)) * input_data) == input_data);
    assign temp_1 = ((input_data ^ input_data) | (~temp_0));
    assign temp_2 = ((temp_0 | input_data) + temp_0);
    assign temp_3 = ((temp_1 | temp_0) ^ temp_1);
    assign temp_4 = (((temp_2 * temp_2) * temp_3) * input_data[3:3]);
    assign temp_5 = ((((temp_1 + temp_2) - (~temp_1)) | input_data) ^ temp_4);
    assign temp_6 = $signed((((temp_1[20:0] << temp_5) | (~temp_1)) & temp_5));
    assign temp_7 = (temp_4 | temp_6);
    assign temp_8 = ((((((temp_6[9:0] & temp_6) * (~temp_0)) <= temp_2) ^ temp_5) - temp_0) + temp_6);
    assign temp_9 = temp_4 ? (((temp_5 | temp_1) << (~temp_5)) * temp_6[3:0]) : ((temp_7 | temp_0) - (~temp_0));
    assign temp_10 = (((((temp_6 + temp_3) ^ temp_9) - temp_7) ^ temp_2) - temp_8);

    assign output_data = (temp_6 - temp_5);

endmodule