module top (
    input [11:0] input_data,
    output [8:0] output_data
);

    logic [22:0] temp_0;
    logic [1:0] temp_1;
    logic [29:0] temp_2;
    logic [15:0] temp_3;
    logic [3:0] temp_4;
    logic [10:0] temp_5;
    logic [7:0] temp_6;
    logic [23:0] temp_7;
    logic [30:0] temp_8;
    logic [15:0] temp_9;
    logic [24:0] temp_10;
    logic [6:0] temp_11;
    logic [15:0] temp_12;
    logic [0:0] temp_13;

    assign temp_0 = ($signed(input_data) + input_data);
    assign temp_1 = temp_0;
    assign temp_2 = temp_0;
    assign temp_3 = temp_1;
    assign temp_4 = ($unsigned(($signed(temp_3) + temp_1)) & temp_2);
    assign temp_5 = temp_1;
    assign temp_6 = $unsigned(temp_2);
    assign temp_7 = {13'b0, temp_5};
    assign temp_8 = input_data;
    assign temp_9 = ($signed(input_data) & temp_5);
    assign temp_10 = (temp_8 * temp_5);
    assign temp_11 = ($unsigned((temp_2[29:18] * temp_4)) * temp_5);
    assign temp_12 = $signed(((temp_5 ^ temp_10) ^ temp_4));
    assign temp_13 = temp_7;

    assign output_data = ($signed(temp_7) - temp_9);

endmodule