module top (
    input [2:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;
    logic [1:0] temp_17;

    assign temp_0 = (input_data + input_data);
    assign temp_1 = input_data[2:2] ? $signed((input_data & temp_0)) : ($signed(input_data) + temp_0);
    assign temp_2 = {24'b0, temp_0};
    assign temp_3 = input_data;
    assign temp_4 = ((temp_0 & (~temp_2)) + temp_2);
    assign temp_5 = temp_1;
    assign temp_6 = input_data[1:1] ? ($signed(($signed(temp_3) & temp_3)) - input_data[2:1]) : (input_data[1:0] & temp_3);
    assign temp_7 = (($unsigned(temp_6) & 26'd25670156) * temp_0);
    assign temp_8 = 19'd399596;
    logic [18:0] expr_35843;
    assign expr_35843 = temp_8;
    assign temp_9 = expr_35843[3:0];
    assign temp_10 = temp_2;
    assign temp_11 = ($unsigned(temp_6) & temp_7);
    assign temp_12 = ($signed(($signed(temp_3) & temp_8)) * temp_0[6:3]);
    assign temp_13 = (temp_10[1:0] | temp_8);
    assign temp_14 = (temp_10 | temp_12);
    assign temp_15 = temp_10;
    assign temp_16 = temp_5;
    logic [19:0] expr_139085;
    assign expr_139085 = $unsigned(((temp_12 - temp_14) * temp_8));
    assign temp_17 = temp_3 ? ((temp_12 & temp_9) & temp_12) : expr_139085[1:0];

    assign output_data = $signed(temp_17);

endmodule