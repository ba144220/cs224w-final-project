module top (
    input [2:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;

    assign temp_0 = ($signed((((input_data - input_data) * input_data) * 7'd99)) & input_data);
    assign temp_1 = $signed((((temp_0 + temp_0) ^ temp_0) & (~input_data)));
    assign temp_2 = ($signed(temp_0[6:0]) + input_data);
    assign temp_3 = ((((temp_1 | input_data) * input_data) - temp_0[6:6]) - (~temp_2));
    assign temp_4 = (temp_0 ^ (~input_data));
    assign temp_5 = (((temp_2 & (~input_data)) - input_data) ^ temp_3);
    assign temp_6 = ((temp_4 ^ input_data[2:1]) & (~temp_0[6:5]));
    assign temp_7 = ($signed(((($unsigned(temp_4) > input_data) | temp_1[3:0]) + temp_2[30:18])) | temp_6);
    assign temp_8 = (((((temp_3 & temp_2[30:23]) * (~temp_0[6:3])) ^ temp_1) - input_data) & temp_4);
    assign temp_9 = ((((($unsigned(temp_2) - temp_5) * temp_5) + temp_1) + temp_1) ^ temp_6);

    assign output_data = $unsigned(((((temp_6 * temp_4) & temp_8) - temp_8[12:0]) + temp_4));

endmodule