module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;
    logic [17:0] temp_12;
    logic [2:0] temp_13;
    logic [1:0] temp_14;
    logic [23:0] temp_15;

    assign temp_0 = ((((($signed(input_data) | (~input_data)) | input_data) & input_data) & input_data) | input_data);
    assign temp_1 = $signed(($signed(($signed(($signed(($signed((($signed((temp_0 * input_data)) * input_data) ^ input_data)) - input_data)) + input_data)) & input_data)) + temp_0));
    assign temp_2 = $signed(11'd463);
    assign temp_3 = (($signed(($unsigned(($signed(($unsigned((((input_data & (~input_data)) - temp_1) * temp_1)) * temp_0)) + input_data)) | (~input_data))) & temp_0[5:1]) - temp_2);
    assign temp_4 = ((($signed(($unsigned(($unsigned((temp_3 - temp_3)) | (~input_data))) | temp_0[5:4])) + (~temp_2)) ^ temp_3) - (~temp_2));
    logic [29:0] expr_462614;
    assign expr_462614 = ($unsigned(($unsigned((($signed(($unsigned(($unsigned((temp_2 & input_data)) * temp_1)) | (~input_data))) & input_data) ^ (~input_data))) | input_data)) * temp_1);
    assign temp_5 = expr_462614[13:0];
    assign temp_6 = (($unsigned((($unsigned(($unsigned(((((temp_0 ^ temp_3) ^ input_data) ^ temp_5) & temp_0)) - input_data)) & input_data) ^ temp_0)) + input_data) + temp_2);
    assign temp_7 = $unsigned(($unsigned((input_data + temp_3)) > temp_5));
    assign temp_8 = $signed((((($signed(input_data) & temp_2) - temp_0[5:4]) * temp_7) - input_data));
    assign temp_9 = (($signed((((temp_4 & temp_5) ^ input_data) + temp_6)) + input_data) * temp_6);
    assign temp_10 = $signed(($unsigned(((($unsigned((temp_2 - (~temp_4[16:8]))) * (~temp_9[25:3])) | temp_1) + temp_7)) + (~temp_8)));
    assign temp_11 = $unsigned((($signed(($signed((($unsigned((((($signed(temp_2) ^ temp_1) * input_data) + (~temp_8)) | input_data)) - temp_0[5:1]) ^ temp_9)) ^ temp_1[23:7])) - temp_6) | temp_4));
    assign temp_12 = (($unsigned(($signed(($signed((($unsigned(((($signed(temp_4) + (~temp_3)) == temp_2[10:8]) * (~temp_11))) < temp_0) + temp_5)) & temp_2)) > temp_9)) | temp_5) * (~temp_4));
    assign temp_13 = input_data[2:2] ? ($unsigned((((temp_1 + temp_9[25:20]) ^ temp_4) - temp_3)) ^ (~temp_6)) : $unsigned((($signed((($signed((($signed(temp_6) + temp_1) - temp_1)) + temp_11) - (~temp_8[27:10]))) | temp_10) & temp_8));
    assign temp_14 = $unsigned(($signed((((((($unsigned(($signed(($signed((temp_9[25:11] & (~temp_0))) ^ temp_8)) | (~temp_9))) + (~temp_9)) | (~temp_3[19:1])) * temp_3) - temp_2) | temp_6) & temp_2[10:5])) ^ temp_10));
    assign temp_15 = (($signed((($unsigned(((((($unsigned(temp_0) | temp_4) ^ temp_13) & temp_10) + temp_7) & temp_12)) - temp_10[23:15]) & temp_5)) * (~temp_10)) * temp_5[13:6]);

    assign output_data = (temp_9 + temp_0);

endmodule