module top (
    input [3:0] input_data,
    output [22:0] output_data
);

    logic [1:0] temp_0;
    logic [29:0] temp_1;
    logic [15:0] temp_2;
    logic [3:0] temp_3;
    logic [10:0] temp_4;
    logic [7:0] temp_5;
    logic [23:0] temp_6;
    logic [30:0] temp_7;
    logic [15:0] temp_8;
    logic [24:0] temp_9;
    logic [6:0] temp_10;
    logic [15:0] temp_11;

    assign temp_0 = input_data[2:2] ? $signed(($signed(input_data[1:0]) - input_data[2:1])) : $signed(($unsigned(input_data[3:2]) ^ input_data[3:2]));
    assign temp_1 = {24'b0, ($unsigned(($signed(temp_0[1:0]) * input_data)) + input_data)};
    assign temp_2 = temp_0[1:0] ? ($unsigned(($unsigned(($unsigned(input_data) | (~input_data))) * input_data)) * input_data) : $unsigned(temp_0);
    assign temp_3 = temp_2;
    assign temp_4 = (($signed(temp_3) - input_data) & temp_1[27:0]);
    assign temp_5 = temp_4;
    assign temp_6 = ($signed(($unsigned(temp_3) ^ temp_2)) ^ temp_2);
    assign temp_7 = (input_data | input_data);
    assign temp_8 = $unsigned(($signed(temp_6) ^ temp_0));
    assign temp_9 = $unsigned(($unsigned(temp_2) < temp_6));
    assign temp_10 = $unsigned(($signed(($unsigned(($signed(($unsigned(temp_1) | input_data)) >> (~temp_9))) + temp_5)) << temp_3));
    assign temp_11 = ($signed(($signed(temp_7) + temp_9)) & temp_4);

    assign output_data = ($unsigned(($signed(($unsigned(temp_11[15:3]) * temp_4)) * temp_10)) + temp_10[6:4]);

endmodule