module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [23:0] temp_0;
    logic [17:0] temp_1;
    logic [8:0] temp_2;
    logic [11:0] temp_3;
    logic [0:0] temp_4;
    logic [21:0] temp_5;
    logic [29:0] temp_6;
    logic [5:0] temp_7;
    logic [21:0] temp_8;
    logic [2:0] temp_9;
    logic [24:0] temp_10;
    logic [10:0] temp_11;
    logic [28:0] temp_12;
    logic [27:0] temp_13;

    assign temp_0 = (((input_data != input_data) & input_data) & input_data);
    assign temp_1 = temp_0 ? $signed(($unsigned(input_data) ^ temp_0)) : ($signed(input_data) + temp_0);
    assign temp_2 = ($signed(($unsigned(($signed(($unsigned(($signed((($signed(($signed(temp_0) >= temp_0)) ^ temp_0) - temp_0[18:0])) != input_data)) < (~temp_1))) * temp_0)) < temp_0)) - input_data);
    assign temp_3 = ($signed(($unsigned(temp_2) + temp_0)) + temp_1);
    assign temp_4 = temp_2;
    assign temp_5 = ($unsigned((($unsigned(($signed(($unsigned(($signed(($unsigned(($signed(temp_1) & temp_0)) ^ temp_3)) & temp_0)) & (~temp_3[2:0]))) & temp_3)) - temp_1) + temp_3)) + temp_4);
    assign temp_6 = $signed(($signed(($unsigned(($signed(($signed(($unsigned(($signed((temp_0 + temp_2)) * 30'd530821750)) & temp_0)) - temp_0)) ^ input_data)) ^ temp_1)) - input_data));
    assign temp_7 = $signed(($signed(temp_6) & temp_4));
    assign temp_8 = $signed(($unsigned(($unsigned(temp_0) << input_data)) & temp_2));
    assign temp_9 = (temp_2 - temp_6[18:0]);
    assign temp_10 = temp_6 ? $unsigned(($signed(($signed((25'd16583682 & input_data)) ^ temp_2[4:0])) * temp_0)) : ($unsigned(($signed(($signed(temp_6) | temp_6[13:0])) ^ temp_1)) * temp_3);
    assign temp_11 = (($unsigned(($unsigned(($unsigned(temp_10) ^ temp_8)) + temp_4)) + temp_6) & temp_10);
    assign temp_12 = {3'b0, ($unsigned(((($signed(temp_8) + (~temp_11)) & temp_11) & temp_4)) & (~temp_0))};
    assign temp_13 = $signed(($unsigned((temp_4 - temp_7)) * temp_8));

    assign output_data = ($unsigned(temp_8) & temp_11);

endmodule