module top (
    input [2:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;
    logic [25:0] temp_16;

    assign temp_0 = input_data[0:0] ? ((input_data ^ input_data) + (~input_data)) : $signed((25'd32793875 & input_data));
    assign temp_1 = $unsigned(temp_0);
    logic [25:0] expr_803707;
    assign expr_803707 = (temp_0 & temp_1[7:0]);
    assign temp_2 = input_data[2:2] ? expr_803707[12:0] : $unsigned((input_data << (~input_data)));
    assign temp_3 = ((temp_0[24:1] * temp_2) + temp_1);
    assign temp_4 = $signed((temp_1 & input_data));
    assign temp_5 = $unsigned((((temp_0 + temp_0) & temp_4) | (~temp_4[5:5])));
    assign temp_6 = temp_5;
    assign temp_7 = ((temp_3 | temp_3) ^ input_data);
    assign temp_8 = temp_7 ? (((input_data | temp_6) & temp_3) ^ temp_6) : (((temp_1[6:0] ^ temp_0[24:5]) + input_data) * temp_1);
    logic [12:0] expr_824632;
    assign expr_824632 = temp_2;
    assign temp_9 = expr_824632[1:0];
    assign temp_10 = $signed((input_data + temp_1));
    assign temp_11 = input_data[2:2] ? $signed(((temp_5 & temp_8[9:0]) - temp_4)) : (temp_6[14:0] * temp_4);
    assign temp_12 = (temp_9[1:1] | temp_5);
    assign temp_13 = ((temp_6 + temp_11) | temp_5[8:3]);
    assign temp_14 = $signed(((temp_7 & temp_7) | temp_5));
    logic [26:0] expr_714644;
    assign expr_714644 = ((temp_0[23:0] - temp_0) ^ temp_0);
    assign temp_15 = temp_12[29:13] ? expr_714644[12:0] : temp_12;
    assign temp_16 = $signed((temp_11 + temp_6));

    assign output_data = $unsigned(((temp_12 ^ temp_6[13:0]) & (~temp_4)));

endmodule