module top (
    input [3:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;

    assign temp_0 = ($unsigned(($unsigned(($unsigned(input_data) ^ input_data)) ^ (~input_data))) + input_data);
    assign temp_1 = $signed(input_data);
    assign temp_2 = $signed(($signed(($signed(($unsigned(($unsigned((((($unsigned(($signed((($signed(($signed(temp_1) | temp_1)) | input_data) * (~temp_1))) & temp_0)) * input_data) + temp_1[8:2]) - (~input_data)) + input_data)) * temp_1)) | temp_1)) & (~input_data))) & temp_0));
    assign temp_3 = ((((($signed(($unsigned((((($signed(($signed(temp_1) ^ input_data[2:0])) | temp_0) & temp_1) ^ input_data[3:1]) + temp_1)) & temp_2)) ^ temp_1) * input_data[3:1]) | temp_2) ^ temp_0) + input_data[2:0]);
    assign temp_4 = ($signed(($unsigned(($signed((((((($signed(temp_3) | temp_2) - temp_2[12:4]) * temp_2[12:2]) & (~temp_2[12:12])) - (~temp_1)) ^ temp_1)) & temp_0)) - temp_3)) & temp_2);
    assign temp_5 = ($unsigned(($unsigned(($signed(($unsigned(($unsigned(($signed((temp_4 * input_data)) ^ temp_2[12:6])) + temp_1[8:3])) & temp_4[5:5])) * temp_2)) * (~input_data))) - input_data);
    assign temp_6 = ($unsigned(($unsigned(temp_5) & input_data)) ^ temp_1);
    assign temp_7 = (((($unsigned(($signed((($unsigned(($unsigned(($unsigned(($signed((temp_0 * temp_5)) + (~temp_5))) - temp_5[8:4])) + input_data)) & input_data) ^ temp_4[5:4])) + temp_6)) * temp_2) - temp_6) ^ temp_1[8:6]) | temp_3);
    assign temp_8 = (((($signed(($unsigned(($signed(($unsigned(($signed(($unsigned(input_data) * temp_4)) & temp_5)) ^ temp_6)) - temp_0)) | temp_2)) ^ input_data) - input_data) + temp_7) ^ temp_6);
    assign temp_9 = $signed((((($signed((($signed(($signed(($unsigned(($signed((((temp_8 & temp_4) | temp_6) ^ input_data[2:1])) | (~temp_1))) - (~temp_5))) * temp_8)) * input_data[2:1]) - temp_2)) & (~temp_6)) - temp_3) - temp_8[11:0]) - (~temp_8)));
    assign temp_10 = (temp_4 + temp_4);
    assign temp_11 = {6'b0, temp_8};
    assign temp_12 = ($signed(($signed((($unsigned(($unsigned(($signed(((($signed(($unsigned(($unsigned(temp_1) + temp_0[24:5])) * temp_10)) - temp_4) * temp_4[5:3]) | temp_9)) ^ temp_0)) * temp_4)) | temp_4) ^ temp_2)) | temp_10)) ^ temp_4);
    assign temp_13 = ($unsigned((($signed(($unsigned(($unsigned((($unsigned((($signed(((temp_0 + temp_5) - temp_12)) & temp_11) | temp_10)) - temp_8) + temp_3)) & temp_9)) - (~temp_10))) ^ temp_0) | temp_10)) + temp_5);

    assign output_data = ($signed((temp_7 & temp_10[19:0])) << temp_2);

endmodule