module top (
    input [3:0] input_data,
    output [9:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;
    logic [26:0] temp_10;
    logic [4:0] temp_11;
    logic [15:0] temp_12;
    logic [5:0] temp_13;
    logic [27:0] temp_14;
    logic [3:0] temp_15;
    logic [7:0] temp_16;
    logic [14:0] temp_17;
    logic [3:0] temp_18;

    assign temp_0 = (($unsigned((input_data | input_data)) == input_data) + input_data);
    assign temp_1 = (($signed(4'd15) ^ input_data) * input_data);
    assign temp_2 = (((input_data ^ temp_0) & temp_1) | temp_0);
    assign temp_3 = (($signed(($signed(input_data) ^ temp_1)) ^ temp_1) | temp_0);
    assign temp_4 = ($signed(($signed((temp_3[1:0] - temp_0[25:1])) * temp_0)) * temp_0);
    assign temp_5 = ($signed(input_data) | temp_0);
    assign temp_6 = ($signed(temp_1) ^ input_data);
    assign temp_7 = (($unsigned(input_data[3:1]) + temp_1) + temp_5);
    assign temp_8 = (temp_6 + temp_2[4:4]);
    assign temp_9 = (($signed(temp_1) < input_data) >= temp_8[5:3]);
    assign temp_10 = {23'b0, ($unsigned(temp_7) - temp_7[2:1])};
    assign temp_11 = ($signed(temp_7) - temp_9);
    assign temp_12 = (($signed(temp_7[2:2]) * temp_3) ^ temp_5);
    assign temp_13 = (temp_5 - temp_0);
    assign temp_14 = 28'd21253744;
    assign temp_15 = (temp_4 | temp_11);
    logic [14:0] expr_768690;
    assign expr_768690 = ($signed(temp_5) * (~temp_6));
    assign temp_16 = temp_8[2:0] ? temp_13 : expr_768690[7:0];
    assign temp_17 = ($unsigned(temp_13) & temp_9);
    assign temp_18 = temp_8[5:4];

    assign output_data = (temp_5 | temp_11);

endmodule