module top (
    input [4:0] input_data,
    output [2:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;

    assign temp_0 = input_data;
    assign temp_1 = input_data[3:0];
    assign temp_2 = input_data;
    assign temp_3 = temp_2;
    assign temp_4 = ($signed(($signed(($signed(($signed(($signed(($signed(temp_2) ^ temp_0)) + input_data)) & temp_0)) ^ temp_3)) - temp_3)) & temp_3);
    assign temp_5 = ($signed(($unsigned(($signed(temp_1[3:3]) - temp_0)) | input_data[3:0])) ^ input_data[4:1]);
    assign temp_6 = {10'b0, temp_1};
    assign temp_7 = ($unsigned((($signed(temp_2[4:4]) & temp_2[4:3]) | temp_4)) * input_data[4:2]);
    assign temp_8 = ($signed(($unsigned((($signed(temp_3) ^ temp_3) * temp_5)) * temp_1)) + temp_5[3:3]);

    assign output_data = ($unsigned(($unsigned(($unsigned(($signed(($unsigned(temp_6) + temp_2)) - temp_7)) ^ temp_1)) - temp_0)) & temp_2);

endmodule