module top (
    input [7:0] input_data,
    output [4:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;
    logic [26:0] temp_10;
    logic [4:0] temp_11;
    logic [15:0] temp_12;
    logic [5:0] temp_13;

    assign temp_0 = input_data;
    logic [25:0] expr_598951;
    assign expr_598951 = temp_0;
    assign temp_1 = expr_598951[3:0];
    assign temp_2 = (((((input_data[7:3] == input_data[7:3]) | temp_0) ^ input_data[4:0]) ^ temp_1) ^ temp_1);
    assign temp_3 = input_data[7:1];
    assign temp_4 = {23'b0, (((((temp_0 | (~temp_1)) < temp_1) ^ (~input_data)) & (~24'd6118411)) < temp_2)};
    assign temp_5 = ((((((((temp_3[1:0] - temp_0[25:1]) * temp_0) * temp_3[4:0]) & temp_1[2:0]) ^ temp_0) + input_data[3:0]) * input_data[4:1]) * temp_4);
    assign temp_6 = ((((((((input_data * temp_4) * temp_0) | (~input_data)) ^ (~temp_3)) ^ temp_5) - (~14'd15248)) | input_data) + temp_5);
    assign temp_7 = ((((input_data[6:4] & 3'd7) | (~temp_4[5:0])) & input_data[3:1]) ^ temp_0);
    assign temp_8 = ((((temp_0 > temp_3) & temp_4) < temp_7) | input_data[5:0]);
    assign temp_9 = (((((((temp_7 - temp_6) + temp_0) | (~temp_8[5:2])) * temp_2[4:4]) * (~temp_8)) + temp_2[4:1]) + temp_3[1:0]);
    assign temp_10 = ((input_data + temp_4) == (~temp_5));
    assign temp_11 = (((temp_6 & input_data[5:1]) ^ (~temp_2)) + temp_4[23:22]);
    assign temp_12 = ((((temp_0 <= (~temp_0)) < (~temp_4)) | temp_2[4:1]) - temp_8[5:5]);
    assign temp_13 = ((temp_10 <= (~temp_8)) == (~temp_11));

    assign output_data = (((((((temp_10 * (~temp_0[25:17])) | temp_1) - temp_11) & temp_1) ^ temp_3[2:0]) ^ temp_4[23:16]) ^ temp_1);

endmodule