module top (
    input [2:0] input_data,
    output [2:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;
    logic [17:0] temp_12;
    logic [2:0] temp_13;
    logic [1:0] temp_14;
    logic [23:0] temp_15;

    assign temp_0 = ((((($signed(input_data) | input_data) | input_data) & input_data) & input_data) | input_data);
    assign temp_1 = {13'b0, (($unsigned(((($unsigned(((input_data * input_data) * input_data)) | temp_0) + temp_0) | temp_0)) ^ input_data) + temp_0)};
    assign temp_2 = (((temp_0 | temp_0) >> (~input_data)) * temp_1);
    assign temp_3 = ((temp_0[2:0] | input_data) & temp_0);
    assign temp_4 = temp_0;
    assign temp_5 = ((($signed(((((temp_1 | temp_4[14:0]) + input_data) | temp_2) - (~input_data))) ^ temp_1) ^ temp_3) * temp_0);
    assign temp_6 = (($unsigned((($signed(($signed(($unsigned((temp_2 * temp_4)) & input_data)) ^ input_data)) & input_data) ^ input_data)) | input_data) * temp_1);
    assign temp_7 = ($unsigned(((($signed((((temp_5 & temp_2) | temp_5) | temp_3)) * temp_5) - input_data) | input_data)) + temp_3);
    assign temp_8 = (temp_5 & temp_1);
    assign temp_9 = ((input_data + temp_7) > temp_4);
    assign temp_10 = ((($signed(($signed(($unsigned(temp_6) | temp_6)) + temp_7)) & input_data) & input_data) ^ temp_4);
    assign temp_11 = ((temp_6 * input_data) ^ input_data);
    assign temp_12 = ((((temp_2 + temp_2) & temp_5) ^ input_data) - temp_5);
    assign temp_13 = ((((($unsigned(temp_2) & temp_2) & temp_0) | temp_9) ^ temp_6) | temp_10);
    assign temp_14 = ($unsigned(((temp_1 & temp_7) | temp_0)) ^ temp_3[16:0]);
    assign temp_15 = ((((((temp_14 ^ temp_1) - temp_6) + temp_7) & temp_11) - temp_9[5:0]) ^ temp_8[25:0]);

    assign output_data = ($signed(temp_5) ^ temp_14);

endmodule