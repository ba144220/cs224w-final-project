module top (
    input [3:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;

    assign temp_0 = ((((((input_data & input_data) & input_data) + input_data) + input_data) ^ input_data) + input_data);
    assign temp_1 = ($unsigned((($unsigned(($unsigned((((input_data | input_data) - temp_0) ^ temp_0[24:11])) * temp_0)) - input_data) - temp_0[19:0])) | temp_0[22:0]);
    assign temp_2 = ((((($unsigned((($signed(($unsigned((temp_1 | temp_1[8:0])) + input_data)) - temp_0) >> temp_1)) ^ temp_0) + temp_1) & (~temp_1)) | input_data) << input_data);
    assign temp_3 = (input_data[3:1] - temp_2);
    assign temp_4 = (($unsigned(((((temp_0 ^ input_data) * temp_2) - input_data) | input_data)) ^ temp_3) + temp_3);
    assign temp_5 = $unsigned(($unsigned(($signed(($unsigned(((temp_1 + input_data) * temp_0)) & temp_0[8:0])) - temp_0[24:0])) * input_data));
    assign temp_6 = ($signed((temp_3 & temp_3)) ^ temp_2);
    assign temp_7 = (($unsigned((($signed((((($unsigned(temp_1) - temp_5) * temp_5[3:0]) - temp_1) + temp_4[5:0])) * temp_2) * input_data)) + temp_5) & temp_4);
    assign temp_8 = (((((((temp_7 ^ temp_2) & temp_6) | temp_1) & temp_3[2:2]) * temp_0) + temp_3) + temp_1);
    logic [30:0] expr_803008;
    assign expr_803008 = ((((((($unsigned((temp_3 * temp_5)) + temp_6) & temp_0) - temp_0) & temp_1) | temp_3) * temp_2) + temp_7);
    assign temp_9 = temp_1 ? ($signed((((($unsigned(temp_6) + temp_7) * temp_0) - temp_7) & temp_8)) | input_data[3:2]) : expr_803008[1:0];
    assign temp_10 = ($signed(($signed(($unsigned((((temp_2 | temp_2) | temp_8) * temp_0)) | temp_7)) ^ temp_1)) | temp_3);

    logic [35:0] expr_153875;
    assign expr_153875 = ((((((($signed(temp_1[8:0]) & temp_9) * temp_10) & temp_10) - temp_7) - temp_3[2:2]) - temp_8) - temp_3[2:1]);
    assign output_data = expr_153875[11:0];

endmodule