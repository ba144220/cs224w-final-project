module top (
    input [2:0] input_data,
    output [36:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;

    assign temp_0 = input_data[1:1] ? ((((($signed((((($unsigned(input_data) - (~input_data)) << input_data) >> input_data) >> input_data)) - input_data) << input_data) >> (~input_data)) & input_data) ^ 5'd6) : input_data;
    assign temp_1 = input_data;
    assign temp_2 = ((((input_data | input_data) | temp_1) | input_data) | temp_0);
    assign temp_3 = temp_0 ? ($unsigned(($signed(($unsigned((temp_0 * temp_2)) + temp_1)) & (~input_data))) * temp_2) : {24'b0, $signed(temp_2)};
    assign temp_4 = temp_2 ? (((($unsigned(input_data) >= temp_0) & temp_3) | temp_1) < temp_0) : $signed((($unsigned((($signed((((($unsigned(temp_1) * temp_2) ^ input_data) & input_data) & temp_1)) | input_data) | temp_0)) | temp_0) & input_data));
    assign temp_5 = temp_2 ? ($unsigned(($signed(((((input_data - temp_4) ^ temp_4) - input_data) | temp_1)) ^ temp_4)) - temp_0[4:1]) : (((($unsigned((($signed(($signed((temp_1 - input_data)) | temp_1)) ^ input_data) ^ input_data)) & temp_4) & temp_3[31:23]) - temp_2) + temp_2);
    assign temp_6 = (((((((temp_4 * input_data) * temp_1) ^ temp_3) | temp_1) + temp_3) ^ input_data) * temp_0);
    assign temp_7 = $unsigned(($signed(($signed((temp_3 & temp_3)) + temp_2)) + temp_4));
    assign temp_8 = ((temp_3 * temp_0) ^ input_data);
    assign temp_9 = temp_8;

    assign output_data = ((((((temp_4 ^ temp_8) ^ temp_4) | temp_0) | (~temp_9)) ^ temp_3) ^ temp_2);

endmodule