module top (
    input [3:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;

    assign temp_0 = ($unsigned(($unsigned(($signed(input_data) - input_data)) ^ input_data)) & input_data);
    assign temp_1 = $unsigned(($unsigned(temp_0) & input_data));
    assign temp_2 = ($signed((temp_0 * temp_0)) * temp_0);
    assign temp_3 = $signed(input_data[2:0]);
    assign temp_4 = $unsigned(($signed(($signed(input_data) & temp_0)) * temp_3));
    assign temp_5 = ($signed(($signed(temp_4[5:0]) * temp_3)) * temp_0);
    assign temp_6 = ($signed((temp_0 + temp_3)) & temp_2);
    assign temp_7 = ($signed(((temp_5 * temp_5) + temp_2)) & temp_6);
    assign temp_8 = ($signed(($unsigned(((temp_7 << temp_4) << temp_3)) & temp_1)) + temp_2[4:0]);
    assign temp_9 = 2'd0;
    assign temp_10 = {4'b0, ((temp_0 | temp_5) << (~temp_4))};
    assign temp_11 = ($signed(($signed(temp_8) * temp_5)) - temp_2);

    assign output_data = ($signed((temp_9 * temp_11)) | temp_2);

endmodule