module top (
    input [5:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;

    assign temp_0 = (input_data ^ input_data);
    assign temp_1 = input_data[3:3] ? {3'b0, input_data} : input_data;
    assign temp_2 = $unsigned(((temp_0 * input_data) * temp_0));
    assign temp_3 = input_data[3:1];
    assign temp_4 = input_data[0:0] ? $unsigned((temp_3 << input_data)) : temp_2;
    assign temp_5 = ($unsigned(temp_4) ^ 9'd215);
    assign temp_6 = $signed((temp_0 & input_data));
    assign temp_7 = $unsigned(($signed((($signed(temp_0) + temp_0) + input_data)) & input_data));
    assign temp_8 = temp_5;
    assign temp_9 = $signed(input_data[3:2]);
    assign temp_10 = (((($unsigned(($signed(temp_9) - temp_8)) & temp_9) * input_data) | temp_3) & temp_1);
    assign temp_11 = temp_10 ? (((32'd2803363716 * temp_1) - temp_9) + temp_1) : $unsigned(((((($signed(temp_4) & temp_0[24:0]) | temp_8) * temp_3) >> temp_9) ^ temp_7));
    assign temp_12 = {2'b0, (($signed(temp_8) | (~temp_2)) * temp_4)};
    assign temp_13 = ($signed((($signed((temp_9 + temp_8[20:0])) * temp_5) * (~temp_12))) - temp_10);

    assign output_data = $signed((($unsigned((($unsigned((temp_7 | temp_7)) - temp_7) >> temp_5)) * temp_12) & temp_2));

endmodule