module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;

    assign temp_0 = input_data[2:2] ? input_data : input_data;
    assign temp_1 = ($signed(temp_0) - input_data);
    assign temp_2 = $unsigned(($signed(temp_1) + temp_1));
    assign temp_3 = temp_2;
    assign temp_4 = ($signed(($signed(temp_1) * temp_2)) ^ temp_0);

    assign output_data = temp_0 ? $signed(($unsigned(temp_3) - temp_0)) : temp_3;

endmodule