module top (
    input [5:0] input_data,
    output [9:0] output_data
);

    logic [23:0] temp_0;
    logic [17:0] temp_1;
    logic [8:0] temp_2;
    logic [11:0] temp_3;
    logic [0:0] temp_4;
    logic [21:0] temp_5;
    logic [29:0] temp_6;
    logic [5:0] temp_7;
    logic [21:0] temp_8;
    logic [2:0] temp_9;
    logic [24:0] temp_10;

    assign temp_0 = {15'b0, ($signed(($signed((input_data + input_data)) ^ input_data)) + (~input_data))};
    assign temp_1 = ($signed(($signed((temp_0[23:19] - input_data)) + temp_0)) ^ temp_0);
    logic [27:0] expr_797692;
    assign expr_797692 = $unsigned(($unsigned((($signed((temp_0 ^ temp_0)) - temp_0) * (~temp_0))) & input_data));
    assign temp_2 = expr_797692[8:0];
    assign temp_3 = ($signed(($signed(temp_1) * (~temp_0))) & temp_1[17:12]);
    assign temp_4 = temp_3;
    assign temp_5 = $signed(($signed((($signed((temp_4 + temp_1)) | temp_1) | input_data)) + input_data));
    assign temp_6 = input_data[5:5] ? ($signed(($unsigned(($signed((temp_2 | temp_1)) & temp_0)) & (~temp_3))) & temp_3) : {7'b0, ($signed(temp_5) + temp_4)};
    assign temp_7 = (((($signed(temp_0) * temp_1) * temp_3) + temp_3) & temp_0);
    assign temp_8 = $unsigned(($unsigned(($unsigned(temp_3) - 22'd3228458)) + temp_6));
    assign temp_9 = $unsigned(temp_1);
    assign temp_10 = $unsigned((((temp_8 * temp_6) - temp_0) + temp_2));

    logic [22:0] expr_581858;
    assign expr_581858 = (temp_1 ^ temp_8);
    assign output_data = temp_4 ? expr_581858[9:0] : temp_7;

endmodule