module top (
    input [3:0] input_data,
    output [9:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;
    logic [0:0] temp_13;
    logic [28:0] temp_14;
    logic [17:0] temp_15;
    logic [14:0] temp_16;

    assign temp_0 = (input_data << input_data);
    assign temp_1 = (((((temp_0 | input_data) ^ input_data) - temp_0) - input_data) ^ input_data);
    assign temp_2 = $signed(temp_1);
    assign temp_3 = $signed((($signed(($signed((((((input_data * temp_2) ^ temp_0) * temp_0) + temp_2) ^ temp_2[1:0])) * temp_2[7:0])) - temp_2[3:0]) - temp_2));
    assign temp_4 = (input_data + temp_3[24:0]);
    assign temp_5 = ((((((((((temp_0 * temp_3[10:0]) + temp_0) * temp_4) | temp_4) ^ input_data) * (~temp_0)) - input_data) ^ temp_3) & input_data) - temp_4);
    assign temp_6 = (((((($signed((((temp_4 + temp_3) | temp_3[18:0]) * temp_2)) + input_data) + temp_4) ^ input_data) * temp_5) + input_data) + temp_2);
    assign temp_7 = (((((((temp_2 * temp_6) & input_data) * temp_0) + input_data) + temp_0) - temp_6) - input_data);
    assign temp_8 = $signed((((temp_5 ^ input_data) - temp_3) | temp_7));
    assign temp_9 = $unsigned((((((((((temp_2[7:0] | (~temp_6[3:0])) <= temp_7) == temp_3) == temp_3[3:0]) ^ temp_3) != temp_7) >= temp_2) + temp_6) != input_data));
    assign temp_10 = ((((((($signed(((temp_7 & input_data[2:1]) - temp_7)) + temp_4) + temp_9) - temp_9) - temp_7) - (~temp_1)) * input_data[3:2]) | (~temp_6));
    assign temp_11 = ((((((temp_1 - temp_4) - input_data) * (~temp_7)) & temp_6) ^ temp_3) ^ temp_6);
    assign temp_12 = ((((((temp_4 + temp_1) + temp_11) | temp_8) | temp_7) ^ input_data) | temp_7);
    assign temp_13 = $signed(temp_6);
    assign temp_14 = $unsigned((((((((((temp_9 - temp_2) + temp_11) + input_data) + temp_8) * temp_11[8:0]) & temp_3) & temp_5) + temp_13) - (~temp_13)));
    assign temp_15 = ((temp_0[1:0] <= temp_0) > temp_11);
    assign temp_16 = ((((((((((temp_5 + temp_13) - temp_2) << temp_1) - temp_1[2:0]) << temp_14[17:0]) ^ temp_1) | temp_3) & temp_10) * temp_14) + temp_9);

    assign output_data = (((($signed(temp_10) * temp_10) ^ temp_10) & temp_11) | temp_1[16:0]);

endmodule