module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;
    logic [17:0] temp_12;
    logic [2:0] temp_13;
    logic [1:0] temp_14;
    logic [23:0] temp_15;
    logic [29:0] temp_16;
    logic [20:0] temp_17;
    logic [24:0] temp_18;

    assign temp_0 = ((6'd17 | input_data) & input_data);
    assign temp_1 = ((($signed((($signed((input_data | input_data)) | input_data) ^ input_data)) * input_data) ^ 24'd282589) ^ temp_0);
    assign temp_2 = ($unsigned(($unsigned((input_data ^ (~temp_0))) + temp_0)) + input_data);
    assign temp_3 = $signed(($unsigned(($unsigned(($signed(($unsigned(input_data) | input_data)) + temp_0)) * temp_2)) * temp_0));
    assign temp_4 = temp_1 ? ($signed(($unsigned(($signed(($unsigned(($signed(17'd107145) - temp_0)) | input_data)) ^ input_data)) | input_data)) | temp_2) : {16'b0, ($unsigned(($unsigned((($signed(($unsigned(($signed(($signed(temp_0[1:0]) ^ temp_0)) * input_data)) ^ input_data)) != input_data) > input_data)) | temp_1)) >= input_data)};
    assign temp_5 = input_data[2:2] ? $unsigned(temp_2) : $unsigned(((($unsigned(($unsigned(((input_data > input_data) * temp_0)) + temp_3)) <= temp_0) == temp_0) * 14'd12641));
    assign temp_6 = ($signed((($signed(temp_5) | temp_5) ^ input_data)) & temp_4);
    assign temp_7 = ($unsigned(($signed(input_data) + temp_3)) == (~temp_5[12:0]));
    assign temp_8 = $signed((($signed((($signed(28'd209984069) | temp_2) - temp_0)) * temp_5[8:0]) & input_data));
    assign temp_9 = $signed(($signed(($signed(($signed(($unsigned((temp_4 << input_data)) ^ (~input_data))) | temp_2)) ^ 26'd47080895)) << temp_5));
    assign temp_10 = temp_3 ? $signed(($unsigned(($signed(($unsigned(($signed(($unsigned(temp_3[19:12]) ^ 24'd2115992)) | temp_1)) & input_data)) | temp_7)) + input_data)) : $unsigned(temp_0[1:0]);
    assign temp_11 = $signed(((($unsigned(((($unsigned(($unsigned(temp_2) + temp_0)) & temp_8[4:0]) ^ temp_9) ^ temp_1)) - temp_6[1:0]) | temp_4) ^ temp_8[27:18]));
    assign temp_12 = temp_11[28:25] ? ($unsigned((($unsigned(temp_3) ^ temp_2) - temp_5)) & input_data) : temp_6;
    assign temp_13 = temp_7 ? ($unsigned(($signed((($signed(($signed((temp_7 | temp_1)) | temp_9)) * temp_12) ^ (~temp_7[8:0]))) | temp_3)) * temp_7) : $signed(($signed(($signed(($signed(($signed((temp_3 * temp_2)) & temp_7)) + temp_8[27:23])) * temp_8)) * (~temp_7[3:0])));
    assign temp_14 = $unsigned((temp_0 >> temp_8));
    logic [30:0] expr_244691;
    assign expr_244691 = (($unsigned(($signed(($signed(temp_2[6:0]) & temp_0)) ^ temp_9)) + (~temp_11)) - temp_14);
    assign temp_15 = expr_244691[23:0];
    assign temp_16 = $unsigned(($signed(temp_8) <= temp_12));
    assign temp_17 = (($unsigned(((($unsigned((temp_14 - temp_4[6:0])) | temp_14) ^ (~temp_12[17:10])) | temp_8)) | temp_7) & temp_7);
    assign temp_18 = (($signed(($signed(($signed(($unsigned((temp_11 - temp_5)) & temp_10)) ^ temp_0[5:4])) * temp_12)) & temp_7) ^ temp_0);

    assign output_data = ($unsigned(($unsigned(($unsigned(temp_10) | temp_15)) * temp_5)) & (~temp_7));

endmodule