module top (
    input [5:0] input_data,
    output [34:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;
    logic [14:0] temp_13;
    logic [9:0] temp_14;
    logic [24:0] temp_15;

    assign temp_0 = 9'd275;
    assign temp_1 = ($signed(($signed(($unsigned(temp_0) * temp_0)) & temp_0)) + input_data);
    assign temp_2 = ($unsigned(($signed(($signed((temp_1[3:0] << (~31'd1783258839))) + (~temp_1))) + temp_0)) ^ temp_0);
    assign temp_3 = ($unsigned(($signed((($signed(temp_1) * temp_0) - temp_2)) * temp_0)) * temp_1);
    assign temp_4 = ($unsigned(($unsigned(($unsigned((temp_2 << temp_0[6:0])) & temp_1[21:0])) - temp_1)) - temp_2);
    assign temp_5 = temp_4;
    assign temp_6 = (($unsigned(($unsigned(temp_2) + temp_2[8:0])) - input_data) * temp_0);
    assign temp_7 = ($signed(($signed((temp_0 * (~temp_2))) << temp_2)) + (~temp_6[4:0]));
    assign temp_8 = ($signed(temp_4) * temp_2);
    assign temp_9 = (($unsigned(($unsigned(temp_0) ^ (~temp_6))) << temp_2) | temp_1);
    assign temp_10 = (($unsigned(((temp_2 | temp_1) + temp_1)) + temp_9) + temp_9);
    assign temp_11 = ($signed(($unsigned(temp_6) - input_data)) | temp_2);
    assign temp_12 = ($unsigned(temp_8) ^ temp_4);
    assign temp_13 = (($unsigned((temp_7 ^ temp_9)) + (~temp_11[13:0])) - temp_10);
    assign temp_14 = ($unsigned(temp_4) - (~temp_11));
    assign temp_15 = temp_3;

    assign output_data = ($unsigned(($unsigned(temp_14) + temp_11)) * (~temp_3));

endmodule