module top (
    input [2:0] input_data,
    output [9:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;

    assign temp_0 = ($unsigned(($unsigned(($unsigned(((($signed((($signed(((((input_data & input_data) - (~input_data)) + input_data) - input_data)) & input_data) * input_data)) ^ 5'd18) ^ input_data) - input_data)) | input_data)) - (~input_data))) - input_data);
    assign temp_1 = ($unsigned(($unsigned((($unsigned((((((temp_0 | temp_0) | input_data) ^ (~temp_0)) * input_data) * temp_0[4:2])) - (~input_data)) + temp_0)) + temp_0)) * temp_0[4:0]);
    assign temp_2 = (($signed(($unsigned(($unsigned(($unsigned(($unsigned((($unsigned((temp_1 - temp_1)) | (~temp_0)) * temp_0)) * input_data)) | input_data)) ^ temp_0)) - temp_1)) + temp_1) + input_data);
    assign temp_3 = ($unsigned(temp_2) | temp_1);
    assign temp_4 = (($signed(($unsigned(((((($signed(temp_3) - temp_3[18:0]) * temp_0) + (~temp_0)) - (~temp_3)) + temp_3)) ^ temp_0)) ^ temp_3) & temp_1);
    assign temp_5 = (($unsigned(($signed(temp_2[7:0]) & temp_4)) * temp_4) | temp_1[8:0]);

    assign output_data = temp_0 ? ($signed(((((((temp_0 + temp_4) * temp_2) - temp_1) | temp_5) - temp_2) * temp_0)) & (~temp_4)) : ($unsigned(($signed((($signed((((((temp_4 | temp_2) + temp_1) == temp_5) & temp_5) | temp_5)) ^ temp_1) <= (~temp_2))) - temp_4)) >= temp_5[30:22]);

endmodule