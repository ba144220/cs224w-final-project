module top (
    input [3:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;
    logic [25:0] temp_16;
    logic [5:0] temp_17;
    logic [31:0] temp_18;

    assign temp_0 = input_data;
    assign temp_1 = temp_0;
    assign temp_2 = ($signed(($unsigned(((temp_0 | temp_1) | temp_1)) - temp_1)) ^ temp_1[8:6]);
    assign temp_3 = ($unsigned(($signed((($signed(($signed(temp_0) * temp_1)) & temp_0) | temp_0)) + temp_0)) * temp_1);
    assign temp_4 = ($unsigned(($signed(($signed(temp_3) & temp_3)) | temp_2[12:1])) ^ temp_0);
    assign temp_5 = ($unsigned((((input_data * temp_0) * temp_3) | temp_2)) * temp_4);
    assign temp_6 = ((($signed(($unsigned((temp_3 + temp_0)) | input_data)) ^ temp_2) | temp_1) ^ temp_4);
    assign temp_7 = $unsigned((((temp_4[5:0] * input_data) + input_data) - temp_4));
    assign temp_8 = ($signed(((temp_6[15:9] - temp_2) ^ temp_2)) & temp_1);
    logic [18:0] expr_911152;
    assign expr_911152 = ($signed(($unsigned((temp_6 * temp_7)) * temp_7)) | temp_3);
    assign temp_9 = expr_911152[1:0];
    assign temp_10 = (($unsigned(temp_2[12:3]) & temp_2) * 30'd791819648);
    assign temp_11 = ($unsigned(temp_5) ^ temp_0);
    assign temp_12 = $unsigned(($unsigned(($unsigned((temp_0 | temp_7)) ^ temp_10[29:24])) * temp_6));
    assign temp_13 = (temp_3[2:2] ^ temp_5);
    assign temp_14 = temp_5[8:4] ? temp_3 : temp_11;
    assign temp_15 = ($unsigned((($signed(temp_3) & temp_2) | temp_12)) ^ input_data);
    assign temp_16 = ($unsigned(($unsigned(($signed(($signed(temp_11) & temp_10)) | temp_10)) - temp_12)) & temp_14[31:11]);
    assign temp_17 = ($unsigned((($unsigned(($signed(temp_3[2:2]) * temp_0)) * temp_5) + temp_14)) ^ temp_16);
    logic [33:0] expr_99050;
    assign expr_99050 = ($signed(($unsigned(($unsigned(((temp_17 & temp_9) | temp_12)) ^ temp_15)) ^ temp_2[12:2])) - temp_14);
    assign temp_18 = expr_99050[31:0];

    assign output_data = ($signed(($signed(temp_3) | temp_14)) * temp_16);

endmodule