module top (
    input [5:0] input_data,
    output [23:0] output_data
);

    logic [17:0] temp_0;
    logic [8:0] temp_1;
    logic [11:0] temp_2;
    logic [0:0] temp_3;
    logic [21:0] temp_4;
    logic [29:0] temp_5;
    logic [5:0] temp_6;
    logic [21:0] temp_7;
    logic [2:0] temp_8;
    logic [24:0] temp_9;
    logic [10:0] temp_10;
    logic [28:0] temp_11;
    logic [27:0] temp_12;
    logic [10:0] temp_13;
    logic [10:0] temp_14;
    logic [15:0] temp_15;

    assign temp_0 = input_data[4:4] ? input_data : input_data;
    assign temp_1 = input_data;
    assign temp_2 = (($unsigned(input_data) & temp_0) & temp_1);
    assign temp_3 = temp_2 ? (temp_2 - input_data[2:2]) : ($signed(temp_0) >= input_data[4:4]);
    assign temp_4 = temp_0;
    assign temp_5 = input_data;
    assign temp_6 = input_data;
    assign temp_7 = $unsigned(($unsigned(temp_0) & temp_0));
    assign temp_8 = temp_6 ? ($signed(($unsigned(input_data[2:0]) + temp_2)) + temp_7) : ($signed(($signed(input_data[2:0]) == temp_4)) + temp_0);
    assign temp_9 = $unsigned(temp_6);
    assign temp_10 = temp_7 ? $signed(($unsigned(($signed(temp_0) - input_data)) - temp_3)) : $signed(temp_4);
    assign temp_11 = ((temp_5 + temp_2) << input_data);
    assign temp_12 = ($signed(input_data) * temp_7);
    assign temp_13 = temp_10;
    assign temp_14 = $signed(($unsigned((temp_5 & temp_13)) & temp_4));
    assign temp_15 = $signed(($unsigned(temp_8) * temp_4));

    assign output_data = ($signed(temp_13) * temp_9);

endmodule