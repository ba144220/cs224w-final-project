module top (
    input [4:0] input_data,
    output [9:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;
    logic [0:0] temp_13;
    logic [28:0] temp_14;
    logic [17:0] temp_15;

    assign temp_0 = (($unsigned((input_data + input_data)) & input_data) & input_data);
    assign temp_1 = ($unsigned(input_data) ^ input_data);
    assign temp_2 = ($unsigned(($signed(($unsigned(($signed(($signed(($signed(($signed(($unsigned(temp_1) | input_data)) - temp_1)) | temp_1)) | temp_1)) ^ temp_0)) | temp_1)) | temp_0)) | (~input_data));
    assign temp_3 = ($unsigned(($signed(($signed(($unsigned(temp_1) | temp_0)) - temp_1)) & (~input_data))) * temp_2);
    assign temp_4 = (($signed(($unsigned(($unsigned(($signed(($unsigned(temp_3) - input_data)) & temp_1[2:0])) & temp_0)) - temp_3)) + temp_2) + input_data);
    assign temp_5 = (temp_4 | temp_2);
    assign temp_6 = ($unsigned(temp_1) | temp_3);
    assign temp_7 = input_data[0:0] ? ($signed(($unsigned((($signed(temp_0) & temp_4) - temp_3)) != temp_0)) != temp_3) : ($unsigned(($unsigned(((($signed(($signed((($unsigned(temp_1) - temp_6) - temp_2)) * (~temp_0))) - temp_2[7:1]) * temp_6) | input_data)) * temp_5)) ^ temp_2);
    assign temp_8 = (($unsigned((($signed(($unsigned(($unsigned(($unsigned((temp_4 & input_data)) & input_data)) | temp_5)) | temp_1[16:11])) ^ temp_3) | temp_4)) ^ input_data) * temp_7);
    assign temp_9 = ((($signed(temp_7) * temp_2) + temp_1) ^ temp_1);
    assign temp_10 = ($unsigned(($unsigned(($unsigned(($unsigned(($unsigned(temp_3) & (~input_data[3:2]))) - temp_9)) * temp_3)) - temp_7)) + 2'd0);
    assign temp_11 = ($unsigned(($unsigned(((temp_5[15:0] ^ temp_4) + temp_6)) ^ temp_8)) ^ input_data);
    assign temp_12 = ($signed(($signed(($unsigned(($signed((($signed(input_data) & input_data) ^ temp_6)) | temp_4)) * (~temp_7))) + temp_0)) * temp_3);
    assign temp_13 = ($signed((($unsigned(($unsigned(($signed(($unsigned(($unsigned(($signed(temp_11) ^ temp_3)) & temp_9)) ^ temp_12)) >> temp_11)) >> (~temp_12))) & (~temp_7)) & temp_7)) ^ temp_4);
    assign temp_14 = ($signed((((temp_11 + temp_1) & temp_4) - temp_0[2:0])) | temp_2);
    assign temp_15 = ($unsigned(temp_2) - temp_6);

    assign output_data = ($unsigned(($signed((($unsigned(($unsigned((temp_1 | (~temp_6))) * temp_2)) + temp_1) * temp_1[16:5])) & temp_0)) & temp_1);

endmodule