module top (
    input [3:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;

    assign temp_0 = (input_data ^ input_data);
    assign temp_1 = temp_0;
    assign temp_2 = (temp_0[19:0] & input_data);
    assign temp_3 = $signed(((input_data[2:0] * temp_2) ^ (~temp_1[8:6])));
    assign temp_4 = (((6'd20 | temp_3) < (~temp_3)) - temp_2[9:0]);
    assign temp_5 = ($unsigned((temp_2 ^ input_data)) | temp_2);
    assign temp_6 = (($signed((temp_0 & input_data)) + temp_0) + input_data);
    assign temp_7 = ((temp_3 | temp_5) ^ (~input_data));
    assign temp_8 = ((temp_5 * temp_3) + temp_4);
    assign temp_9 = ((temp_5 | temp_3) & temp_1);
    assign temp_10 = (temp_4[5:5] * temp_1[8:2]);
    assign temp_11 = temp_5[8:2];
    assign temp_12 = (temp_1[4:0] + (~temp_2));
    assign temp_13 = ((temp_1 - temp_2) & temp_7);

    assign output_data = (((temp_12 ^ temp_7) | temp_8) & (~temp_12[16:0]));

endmodule