module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;
    logic [17:0] temp_12;
    logic [2:0] temp_13;
    logic [1:0] temp_14;
    logic [23:0] temp_15;

    assign temp_0 = (($signed(input_data) | (~input_data)) | input_data);
    assign temp_1 = (($signed(input_data) & temp_0) * temp_0);
    assign temp_2 = ((input_data * temp_1) | input_data);
    assign temp_3 = temp_1 ? $signed(temp_0[5:1]) : temp_2;
    assign temp_4 = $unsigned(input_data);
    assign temp_5 = ((temp_4 << (~input_data)) ^ 14'd4179);
    assign temp_6 = $signed((($unsigned(temp_0) ^ temp_0[2:0]) ^ (~input_data)));
    assign temp_7 = (($signed(temp_0) - temp_5[2:0]) - temp_5);
    assign temp_8 = {12'b0, (((temp_6 - temp_7) | (~temp_5)) & temp_0[5:4])};
    assign temp_9 = temp_1 ? temp_5[13:2] : ($signed(($signed(temp_0) + temp_7)) & temp_6);
    assign temp_10 = temp_5;
    assign temp_11 = temp_10;
    assign temp_12 = ((($signed(temp_4[16:8]) & (~temp_5)) | temp_11) ^ temp_6);
    assign temp_13 = $unsigned((temp_6 + temp_8));
    logic [21:0] expr_747334;
    assign expr_747334 = (temp_12 & temp_9[20:0]);
    assign temp_14 = expr_747334[1:0];
    assign temp_15 = temp_10;

    logic [30:0] expr_584498;
    assign expr_584498 = ((temp_14[1:0] | temp_11) ^ temp_4[16:0]);
    assign output_data = expr_584498[5:0];

endmodule