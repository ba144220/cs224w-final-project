module top (
    input [2:0] input_data,
    output [9:0] output_data
);

    logic [23:0] temp_0;
    logic [17:0] temp_1;
    logic [8:0] temp_2;
    logic [11:0] temp_3;
    logic [0:0] temp_4;
    logic [21:0] temp_5;
    logic [29:0] temp_6;
    logic [5:0] temp_7;

    assign temp_0 = {21'b0, $signed(input_data)};
    assign temp_1 = (input_data - input_data);
    assign temp_2 = input_data;
    assign temp_3 = $signed(($unsigned(input_data) ^ temp_0));
    assign temp_4 = ($unsigned(($signed(input_data[2:2]) ^ temp_1)) & input_data[2:2]);
    assign temp_5 = $signed(($unsigned((($signed((($signed(temp_1) >= temp_3) ^ (~temp_2))) <= temp_3) - input_data)) * temp_1));
    assign temp_6 = $signed(temp_4);
    assign temp_7 = (($unsigned((($signed(temp_5) * (~temp_2)) * temp_5)) & temp_3) | temp_5[19:0]);

    assign output_data = $unsigned(($signed(temp_4) - temp_1[16:0]));

endmodule