module top (
    input [3:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;
    logic [25:0] temp_16;
    logic [5:0] temp_17;

    assign temp_0 = input_data;
    assign temp_1 = $unsigned((temp_0 & input_data));
    assign temp_2 = $signed((((((((((temp_1 - input_data) & temp_0) | (~input_data)) * temp_0) - temp_0) - temp_0) - (~temp_1[8:2])) + temp_1) | temp_0));
    assign temp_3 = $signed((((((((temp_2 & temp_0) & temp_2) + input_data[3:1]) + temp_1) + temp_1) ^ temp_2) + temp_1));
    assign temp_4 = $unsigned((((((temp_2 * temp_0) * temp_3) ^ temp_2) + temp_0) | input_data));
    assign temp_5 = $signed((((input_data * temp_0) & input_data) * temp_3));
    assign temp_6 = temp_2[12:4];
    assign temp_7 = ((((temp_0 & (~temp_2[12:12])) - (~temp_1)) ^ temp_1) & temp_5);
    assign temp_8 = $signed((((((((temp_4 | temp_5) | temp_4) & temp_4) & temp_1[8:6]) & temp_2[12:3]) & temp_1) * input_data));
    assign temp_9 = (((((temp_0 ^ input_data[1:0]) & temp_8[25:9]) ^ temp_4) ^ temp_7) + temp_7);
    assign temp_10 = temp_3;
    assign temp_11 = temp_5[1:0];
    assign temp_12 = $signed(((((((((((temp_5 + temp_10) << input_data) ^ input_data) & input_data) + (~temp_11)) & temp_11[31:26]) >> temp_5) >> input_data) >> temp_8) & temp_10));
    assign temp_13 = $signed((((temp_5 + temp_10) & temp_11) ^ (~temp_8)));
    assign temp_14 = temp_5;
    assign temp_15 = (((((((((((input_data & temp_3) | temp_10) - input_data) | temp_6) * temp_0) | temp_11) + temp_10[29:13]) - temp_5) + temp_4) & temp_4[5:2]) & temp_13);
    assign temp_16 = (temp_13 ^ temp_14);
    assign temp_17 = $unsigned((((((temp_16 & (~temp_9)) - temp_5) + temp_9) & temp_9[1:1]) * temp_13[9:0]));

    assign output_data = temp_3;

endmodule