module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;

    assign temp_0 = input_data;
    assign temp_1 = $signed((input_data & temp_0));
    assign temp_2 = ((temp_1 + temp_1) * temp_0);
    assign temp_3 = ($signed(($signed(temp_0) | temp_0)) + input_data);
    logic [11:0] expr_57955;
    assign expr_57955 = (($signed(temp_3) | input_data) * input_data);
    assign temp_4 = expr_57955[5:0];
    assign temp_5 = ((temp_3 + temp_4) - temp_3);
    assign temp_6 = temp_1;
    assign temp_7 = {22'b0, input_data};
    assign temp_8 = ($unsigned((temp_7 & temp_4)) * input_data);
    assign temp_9 = ((temp_6[1:1] + temp_4) | temp_3);
    assign temp_10 = temp_4;
    assign temp_11 = temp_8;
    assign temp_12 = {17'b0, (temp_5 != temp_1)};
    assign temp_13 = ($unsigned(temp_7) + temp_0);
    assign temp_14 = (temp_10[1:0] | temp_8);

    assign output_data = (temp_9 - temp_6);

endmodule