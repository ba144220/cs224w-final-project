module top (
    input [4:0] input_data,
    output [2:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;

    assign temp_0 = $unsigned(($unsigned(($signed(($signed(input_data) - input_data)) + input_data)) * input_data));
    assign temp_1 = $signed(($unsigned(($signed(($unsigned(((($signed(($unsigned(temp_0) - input_data[4:1])) * input_data[4:1]) & temp_0) ^ temp_0)) & input_data[4:1])) * input_data[4:1])) + temp_0[25:8]));
    assign temp_2 = $signed((($signed(($signed((($signed(($unsigned(temp_1) - temp_0)) * temp_1) | input_data)) ^ input_data)) - temp_0[25:20]) + input_data));
    assign temp_3 = $unsigned((input_data + temp_2));
    assign temp_4 = (($signed((($signed(($signed(($unsigned(($signed(($unsigned(temp_0) * input_data)) - temp_1)) * temp_0)) ^ input_data)) * temp_0) & input_data)) ^ temp_3) + temp_3);
    assign temp_5 = (($signed(temp_0) < input_data[3:0]) >= temp_4);
    assign temp_6 = $unsigned(($signed((($unsigned(($unsigned(($signed(($unsigned(temp_1[3:2]) - temp_1)) | temp_3[6:5])) + temp_4[3:0])) | temp_2) * input_data)) + temp_2[2:0]));
    assign temp_7 = $unsigned(($signed(($signed(($unsigned(($unsigned(($signed(input_data[2:0]) & temp_1)) * temp_2)) + temp_4)) + temp_2[2:0])) ^ temp_2));
    assign temp_8 = $unsigned(($signed(($signed(($signed((temp_1 * temp_7[2:0])) - temp_3)) ^ (~temp_3))) * temp_0));
    assign temp_9 = ($unsigned(($signed(($signed(($unsigned(((($signed(($signed(($signed(($signed(($signed((($signed(temp_3) ^ temp_2) ^ temp_6[13:7])) * temp_4[6:0])) * temp_8[5:3])) + temp_8)) - temp_0)) - temp_6) - temp_8) | temp_0)) ^ temp_1[1:0])) & temp_0)) ^ temp_8)) * temp_3);

    assign output_data = temp_3[2:0] ? (($unsigned(($unsigned(($unsigned(($signed(temp_4) & temp_0)) ^ temp_8)) * temp_1[3:2])) * temp_6) | temp_4) : (($unsigned(($signed(temp_6[1:0]) & temp_7)) * temp_0) + temp_4[23:13]);

endmodule