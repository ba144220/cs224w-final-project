module top (
    input [11:0] input_data,
    output [8:0] output_data
);

    logic [22:0] temp_0;
    logic [1:0] temp_1;
    logic [29:0] temp_2;
    logic [15:0] temp_3;
    logic [3:0] temp_4;
    logic [10:0] temp_5;
    logic [7:0] temp_6;
    logic [23:0] temp_7;
    logic [30:0] temp_8;
    logic [15:0] temp_9;
    logic [24:0] temp_10;
    logic [6:0] temp_11;

    assign temp_0 = $unsigned(input_data);
    assign temp_1 = ($signed(($unsigned(temp_0) - temp_0)) & temp_0);
    assign temp_2 = (temp_1 - temp_0);
    assign temp_3 = ($signed(((($signed((($unsigned((input_data & temp_1)) * 16'd11951) - temp_2)) + temp_2) | 16'd45066) & temp_2[16:0])) ^ temp_0);
    assign temp_4 = $unsigned((((((((($signed((temp_3 * temp_3[15:14])) ^ input_data[5:2]) | temp_2) ^ temp_3) * temp_0) * input_data[8:5]) ^ input_data[5:2]) * input_data[11:8]) * input_data[4:1]));
    assign temp_5 = ($signed((((((input_data[10:0] - temp_3) ^ temp_3) - temp_4[2:0]) + temp_1) & input_data[11:1])) * temp_4);
    assign temp_6 = ($unsigned(((((($signed(($unsigned(temp_1) * input_data[10:3])) - temp_4) & temp_1) & temp_2) | input_data[7:0]) + temp_4)) * input_data[9:2]);
    assign temp_7 = (temp_5 <= (~temp_2));
    assign temp_8 = ((($signed((($unsigned(($signed(($signed((((temp_6 >> temp_6) >> temp_1[1:1]) >> input_data)) ^ temp_6)) - temp_0)) - temp_3) >> (~temp_2))) - temp_1) + temp_5) + temp_4);
    assign temp_9 = (($signed((((((($unsigned(temp_2) & temp_2[29:11]) + temp_7) | temp_6[2:0]) - temp_1) | temp_3) & temp_5)) | temp_3) + temp_7);
    assign temp_10 = ($signed(($unsigned((($signed((((temp_5 >> temp_4[1:0]) + (~temp_0)) + temp_7)) >> temp_2[23:0]) << temp_5)) >> temp_3)) | temp_0);
    assign temp_11 = ((($signed(((($signed((((((temp_7[8:0] ^ temp_6[7:7]) + temp_3) + temp_1[1:0]) - temp_7) ^ temp_0)) - temp_2[29:25]) | temp_3) * temp_3[4:0])) + temp_5) - (~temp_7)) + temp_4[2:0]);

    assign output_data = (((($unsigned((temp_11[6:1] * (~temp_5))) << temp_2) - temp_4) << temp_6[3:0]) << temp_2);

endmodule