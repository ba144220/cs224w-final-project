module top (
    input [2:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;
    logic [12:0] temp_15;
    logic [25:0] temp_16;
    logic [5:0] temp_17;

    assign temp_0 = input_data;
    assign temp_1 = input_data[1:1] ? input_data : input_data;
    assign temp_2 = ($signed(($signed(temp_0) * input_data)) ^ temp_0);
    logic [26:0] expr_147210;
    assign expr_147210 = (($signed(($signed(temp_2[12:3]) * temp_1)) & temp_0) | temp_0);
    assign temp_3 = expr_147210[2:0];
    assign temp_4 = ($unsigned(($signed(($signed(($signed((temp_2[8:0] - temp_0)) - temp_3[2:1])) + temp_3)) | temp_2[12:1])) ^ temp_0);
    assign temp_5 = ($unsigned((((input_data * temp_0) * temp_3) | temp_2)) * temp_4);
    assign temp_6 = ((($signed(($unsigned((temp_3 + temp_0)) | input_data)) ^ temp_2) | temp_1) ^ temp_4);
    assign temp_7 = temp_6 ? ($unsigned(($signed(($unsigned((input_data + input_data)) + input_data)) + temp_0)) - temp_6) : input_data;
    assign temp_8 = input_data;
    assign temp_9 = temp_7 ? ($signed(($signed(($unsigned((input_data[2:1] ^ temp_7)) * temp_7)) | temp_3)) * temp_0) : temp_2;
    assign temp_10 = (($unsigned(temp_5) * temp_7) & temp_0);
    assign temp_11 = $unsigned(($unsigned(($unsigned(($unsigned(temp_10[29:15]) ^ temp_10)) ^ temp_10[29:24])) * temp_6));
    assign temp_12 = ($signed(input_data) + temp_11);
    assign temp_13 = temp_6;
    assign temp_14 = (temp_6 - temp_10);
    assign temp_15 = ($unsigned(($signed(($signed((($unsigned(temp_12) - temp_13) - temp_11)) & temp_13)) | temp_14)) + temp_12);
    assign temp_16 = ($signed(temp_4) & temp_10);
    assign temp_17 = (($unsigned((temp_6[1:0] ^ temp_16)) - temp_14) * temp_10);

    assign output_data = temp_7;

endmodule