module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;

    assign temp_0 = ($signed(($signed(input_data) != input_data)) + input_data);
    assign temp_1 = temp_0;
    assign temp_2 = (($signed(temp_1) & temp_1) | temp_1);
    assign temp_3 = $unsigned(($unsigned(($unsigned(temp_0) & temp_2)) ^ temp_2));
    assign temp_4 = ($signed(($signed(temp_0[5:3]) - temp_0)) ^ temp_0[5:1]);

    assign output_data = temp_4 ? temp_4 : ($signed(temp_0) | temp_1);

endmodule