module top (
    input [4:0] input_data,
    output [36:0] output_data
);

    logic [4:0] temp_0;
    logic [16:0] temp_1;
    logic [7:0] temp_2;
    logic [31:0] temp_3;
    logic [28:0] temp_4;
    logic [30:0] temp_5;
    logic [24:0] temp_6;
    logic [13:0] temp_7;
    logic [6:0] temp_8;
    logic [31:0] temp_9;
    logic [1:0] temp_10;
    logic [24:0] temp_11;
    logic [27:0] temp_12;

    assign temp_0 = ($unsigned(($signed(($unsigned(($signed(($unsigned(($signed(input_data) | input_data)) & input_data)) & input_data)) * input_data)) - input_data)) ^ input_data);
    assign temp_1 = ($signed(($signed(($signed(($unsigned(temp_0) | (~input_data))) - temp_0)) | temp_0)) | temp_0);
    assign temp_2 = ($signed(($unsigned(($unsigned(($signed(($unsigned(($signed(temp_0) & input_data)) & input_data)) & temp_0)) * temp_0[1:0])) * temp_0[4:2])) ^ input_data);
    assign temp_3 = ($unsigned(($unsigned(temp_2) - temp_0[2:0])) - input_data);
    assign temp_4 = temp_0;
    logic [31:0] expr_450091;
    assign expr_450091 = ($unsigned(($unsigned(($signed(temp_0) | temp_4)) & (~temp_3[22:0]))) | input_data);
    assign temp_5 = expr_450091[30:0];
    logic [35:0] expr_702977;
    assign expr_702977 = ($signed(($unsigned(($signed(($unsigned(($unsigned(temp_5) | temp_5[5:0])) * temp_2)) ^ input_data)) - input_data)) * temp_2);
    assign temp_6 = expr_702977[24:0];
    logic [19:0] expr_332765;
    assign expr_332765 = ($signed(($signed(($signed(temp_1) - temp_1)) | input_data)) * temp_0);
    assign temp_7 = expr_332765[13:0];
    logic [33:0] expr_577980;
    assign expr_577980 = ($signed(($signed(($unsigned(temp_7) | (~temp_3[31:9]))) | temp_3)) * (~temp_1));
    assign temp_8 = expr_577980[6:0];
    assign temp_9 = ($unsigned(($unsigned(($unsigned(($signed(($unsigned(temp_5) - temp_5[22:0])) * temp_8)) ^ temp_5)) ^ temp_4)) + temp_7);
    assign temp_10 = 2'd1;
    assign temp_11 = $unsigned(($signed(($signed(($unsigned(($unsigned((($signed(temp_1[16:11]) | temp_7) - temp_5)) ^ temp_1)) - temp_4)) + temp_8)) + temp_6));
    assign temp_12 = $signed(($unsigned(($signed(temp_9) - temp_3)) ^ temp_9));

    assign output_data = temp_9[21:0];

endmodule