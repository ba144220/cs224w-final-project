module top (
    input [2:0] input_data,
    output [17:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;
    logic [14:0] temp_13;
    logic [9:0] temp_14;
    logic [24:0] temp_15;
    logic [0:0] temp_16;

    assign temp_0 = (input_data * input_data);
    assign temp_1 = $unsigned(((temp_0 | temp_0) ^ input_data));
    assign temp_2 = ((($signed(((($signed((($unsigned(($unsigned(input_data) * temp_1)) - (~temp_1)) ^ input_data)) * temp_0) - input_data) & temp_1)) | temp_0) & input_data) + input_data);
    assign temp_3 = temp_2[12:0] ? ($unsigned(($unsigned(((input_data * input_data) + input_data)) * temp_0)) ^ input_data) : ($unsigned(temp_2) ^ temp_2);
    assign temp_4 = $unsigned(((((((temp_3 | temp_1[15:0]) | input_data[0:0]) * temp_1[23:0]) & temp_0) + temp_3[1:0]) | temp_0));
    assign temp_5 = temp_2;
    assign temp_6 = temp_0 ? input_data : ((temp_4 * (~temp_1)) - temp_3);
    assign temp_7 = ($unsigned(($signed(($unsigned(($unsigned((($unsigned((input_data - temp_2)) + input_data) ^ temp_4)) + (~input_data))) + temp_5)) + temp_6)) | temp_5);
    assign temp_8 = input_data[1:1] ? ((($unsigned(((((((temp_6 + temp_3) ^ temp_7) & input_data) - temp_3) | input_data) * input_data)) - temp_3) | temp_0) ^ input_data) : $unsigned(((($signed(temp_4) ^ input_data) + (~temp_1)) & temp_5[11:0]));
    assign temp_9 = ((temp_6 * temp_5) ^ temp_4);
    assign temp_10 = $signed(temp_2);
    assign temp_11 = ($signed((((($unsigned(((temp_5 & temp_10) + temp_8)) & temp_2[17:0]) * input_data) + temp_9) - temp_9)) | temp_6);
    assign temp_12 = ($signed(((($unsigned(($unsigned(((temp_8 & input_data) + temp_11)) - temp_7)) & temp_4) + temp_9) * temp_5)) + temp_11);
    assign temp_13 = temp_6;
    assign temp_14 = (($signed(((temp_7 ^ temp_13) + temp_4)) - temp_9) & (~temp_13[8:0]));
    assign temp_15 = temp_14 ? (temp_1 + temp_4) : (($unsigned(($unsigned(temp_5) << (~input_data))) + temp_3) >> temp_10[10:0]);
    assign temp_16 = ((((((temp_12 ^ temp_11) ^ temp_8) ^ (~temp_15[6:0])) & (~temp_3)) | temp_14) + temp_12);

    assign output_data = $unsigned(temp_4);

endmodule