module top (
    input [3:0] input_data,
    output [9:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;
    logic [26:0] temp_10;
    logic [4:0] temp_11;

    assign temp_0 = ($signed(((((($unsigned(((input_data ^ input_data) - input_data)) + input_data) + input_data) & input_data) & input_data) - input_data)) ^ input_data);
    assign temp_1 = temp_0 ? (($signed((($signed((((input_data ^ temp_0) & temp_0) | temp_0)) & temp_0) ^ (~temp_0))) - temp_0[19:0]) | temp_0) : (((((((($unsigned((((((temp_0 & (~temp_0)) | temp_0) + input_data) | temp_0) * temp_0)) | temp_0) + temp_0) | temp_0) - temp_0) + input_data) * temp_0) - temp_0) ^ temp_0);
    assign temp_2 = (((($signed((((($unsigned(((input_data ^ (~input_data)) | input_data)) & temp_1) + temp_0) * temp_0) + input_data)) | temp_0) + temp_0) * temp_1) * temp_0);
    assign temp_3 = ((((((((temp_1 | input_data) - temp_0) & temp_2) ^ temp_0) + temp_1) | (~temp_1)) | temp_2[3:0]) + (~temp_0));
    assign temp_4 = $unsigned(($signed((($unsigned((($unsigned((input_data ^ (~temp_2[2:0]))) + temp_2[2:0]) * (~input_data))) ^ temp_0) | temp_2)) * temp_0));
    assign temp_5 = ($unsigned(((((((((($unsigned(($signed((($signed(temp_1) ^ (~temp_1)) ^ temp_3[6:4])) * temp_2[2:0])) * input_data) - temp_3[3:0]) | temp_0[25:13]) * temp_1[3:0]) ^ temp_4) ^ temp_1[3:0]) ^ temp_4) + temp_4) + temp_1)) + temp_4);
    assign temp_6 = (temp_2 - temp_3);
    assign temp_7 = (temp_5 + temp_3);
    assign temp_8 = $unsigned((($unsigned((((($unsigned((temp_4 + temp_1)) - temp_3[1:0]) - temp_4) & temp_2[4:0]) ^ temp_5)) * temp_1) + (~temp_1)));
    assign temp_9 = (((temp_5 + temp_6) + temp_6) + temp_8);
    assign temp_10 = (($signed(((((((((temp_1 - temp_7) & temp_3) * temp_9[27:14]) - temp_5) ^ temp_3[2:0]) & temp_0) | temp_1) & (~temp_1))) ^ temp_7[1:0]) + temp_4);
    assign temp_11 = $unsigned(($unsigned((($signed(((((($signed((temp_0[10:0] & temp_5)) - temp_6) & (~temp_3)) * temp_5) | temp_7) - temp_4[20:0])) - temp_10[20:0]) | temp_0)) * temp_1));

    assign output_data = (((($unsigned((temp_1 + temp_8)) & temp_1[2:0]) * temp_5) ^ temp_6[1:0]) + temp_4[23:20]);

endmodule