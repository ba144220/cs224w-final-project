module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;
    logic [1:0] temp_17;
    logic [16:0] temp_18;

    assign temp_0 = (input_data + input_data);
    assign temp_1 = ($unsigned(($signed((($unsigned(temp_0) << (~temp_0)) + temp_0)) & temp_0)) & 26'd30718336);
    assign temp_2 = $signed(input_data);
    assign temp_3 = (($signed((10'd909 * temp_1)) & temp_1) + temp_0);
    assign temp_4 = input_data;
    assign temp_5 = {1'b0, input_data};
    assign temp_6 = (temp_2[2:0] * temp_4);
    assign temp_7 = ($unsigned(input_data) ^ temp_5);
    assign temp_8 = ((temp_2 + input_data) & temp_0);
    assign temp_9 = ($unsigned(temp_5) & input_data);
    assign temp_10 = ($unsigned((input_data - temp_8)) > input_data);
    assign temp_11 = {23'b0, ($signed(($signed(($signed(temp_4) - input_data)) ^ temp_0[6:3])) >= temp_1)};
    assign temp_12 = ((temp_9 & temp_7) * temp_1);
    assign temp_13 = (((((temp_2 * (~temp_0)) ^ temp_1[19:0]) - temp_1[16:0]) | temp_11) | temp_11);
    assign temp_14 = ($unsigned(($unsigned(temp_8) * temp_6)) * temp_4);
    assign temp_15 = temp_12;
    assign temp_16 = temp_3 ? input_data : ($signed(temp_0) | temp_6);
    assign temp_17 = (($unsigned((temp_0 * temp_4[1:0])) - temp_0) ^ temp_12);
    assign temp_18 = (((((temp_6 ^ temp_15) * temp_1) + temp_1) - temp_10) | (~temp_2));

    assign output_data = ($signed(temp_11) & temp_12[14:0]);

endmodule