module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;
    logic [17:0] temp_12;
    logic [2:0] temp_13;

    assign temp_0 = ((((($signed(input_data) | input_data) | input_data) & input_data) & input_data) | input_data);
    assign temp_1 = $unsigned(((((($unsigned(((input_data * input_data) * input_data)) | temp_0) + temp_0) | temp_0) ^ (~24'd8371887)) + temp_0[5:2]));
    assign temp_2 = $signed(input_data);
    assign temp_3 = ((((($unsigned(((((((temp_2 & temp_2[10:8]) <= temp_1) | temp_1) | temp_0) != (~input_data)) - temp_2)) | (~temp_0)) - temp_0[5:1]) | temp_1) < temp_0[5:4]) - input_data);
    assign temp_4 = $signed((((((temp_0 ^ input_data) - input_data) ^ temp_3) * temp_0[5:5]) - 17'd11319));
    assign temp_5 = $unsigned((((($unsigned((($signed(($signed((input_data ^ temp_1)) ^ input_data)) & input_data) ^ input_data)) | input_data) * temp_1) | input_data) ^ temp_4));
    assign temp_6 = $unsigned((((($signed((($unsigned(($unsigned(((($signed((input_data | temp_3)) * temp_5) - temp_4) | input_data)) + temp_3)) + temp_3) * temp_4)) & temp_5) & (~temp_1[18:0])) + temp_3) - temp_4));
    assign temp_7 = $signed((((($signed((((($unsigned(temp_3) - input_data) | temp_0) * temp_2) - input_data)) + input_data) * input_data) * input_data) ^ input_data));
    assign temp_8 = $signed((((((input_data * input_data) << temp_5) * temp_3[19:5]) * temp_4) + temp_5));
    assign temp_9 = (((((((($signed(($unsigned(temp_6[2:2]) & temp_5)) & input_data) + temp_2) & (~temp_0)) & temp_1) & (~temp_7[10:9])) | input_data) - temp_0[5:1]) | temp_6);
    assign temp_10 = $signed((($unsigned((($signed(((((temp_3 ^ temp_6) - temp_4) * temp_1) >= temp_2)) + temp_3) == temp_2[10:8])) * temp_4) + (~temp_1)));
    logic [34:0] expr_406052;
    assign expr_406052 = ((($unsigned(((((($unsigned(($unsigned(($signed((temp_2 & input_data)) & temp_7)) & temp_9)) | (~temp_4)) | temp_10) + temp_9[25:20]) ^ temp_4) - temp_3)) ^ temp_6) | temp_6) * temp_3);
    assign temp_11 = expr_406052[28:0];
    assign temp_12 = $unsigned(($signed(((((($signed(temp_5) | temp_7) - temp_3) + temp_8) * temp_4) + temp_1)) * temp_4));
    assign temp_13 = $unsigned((((((((($unsigned(((temp_6 * temp_0[3:0]) + temp_9)) - (~temp_1)) | temp_3) * temp_2) <= temp_6) > temp_2[10:5]) == temp_10) | temp_5) + temp_0));

    assign output_data = ($signed(((((((temp_13 * temp_6) ^ temp_6) ^ temp_13) * temp_12) - temp_6) * temp_5)) * temp_10[23:19]);

endmodule