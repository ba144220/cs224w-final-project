module top (
    input [11:0] input_data,
    output [4:0] output_data
);

    logic [22:0] temp_0;
    logic [1:0] temp_1;
    logic [29:0] temp_2;
    logic [15:0] temp_3;
    logic [3:0] temp_4;
    logic [10:0] temp_5;
    logic [7:0] temp_6;
    logic [23:0] temp_7;

    assign temp_0 = $signed((((input_data & input_data) - (~input_data)) + input_data));
    logic [25:0] expr_786217;
    assign expr_786217 = (((temp_0 - input_data[6:5]) + input_data[2:1]) & (~input_data[8:7]));
    assign temp_1 = expr_786217[1:0];
    assign temp_2 = $signed(((((((temp_0 >= input_data) ^ temp_1) | temp_0) | input_data) - input_data) + temp_1[1:0]));
    assign temp_3 = temp_0[19:0] ? ((temp_1[1:1] * temp_2) ^ temp_1) : (((((((temp_2 * temp_1) ^ temp_1) * temp_2) * temp_2) ^ input_data) * input_data) & temp_0);
    assign temp_4 = $unsigned(((((((((temp_0 | temp_1) - temp_1[1:0]) & temp_3) * temp_3) | temp_0) | temp_2) * temp_1) | temp_0));
    assign temp_5 = ($unsigned(((temp_3 | temp_2) & input_data[10:0])) & temp_0);
    assign temp_6 = ((((temp_3 ^ temp_5[10:3]) * temp_5) | temp_0) | temp_3);
    assign temp_7 = ((($signed((((temp_2 * temp_5) * temp_3) & temp_6[6:0])) + temp_0) + temp_1) * temp_3);

    assign output_data = temp_6 ? (temp_2[3:0] * (~temp_7)) : ((((((((temp_3 * temp_4) ^ (~temp_6)) ^ temp_0[4:0]) & (~temp_7)) ^ temp_6[2:0]) - temp_1[1:0]) | temp_6) * temp_6);

endmodule