module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;
    logic [17:0] temp_12;
    logic [2:0] temp_13;
    logic [1:0] temp_14;
    logic [23:0] temp_15;
    logic [29:0] temp_16;
    logic [20:0] temp_17;

    assign temp_0 = ((($unsigned(input_data) - input_data) | input_data) & input_data);
    assign temp_1 = ($unsigned(input_data) & temp_0);
    assign temp_2 = ($signed(($signed((((input_data | temp_1) | temp_1) | input_data)) - input_data)) + input_data);
    assign temp_3 = $signed((($unsigned(temp_0[5:1]) * temp_0) - temp_0[5:0]));
    assign temp_4 = ((((input_data & (~input_data)) - temp_3) * input_data) ^ temp_0);
    assign temp_5 = ($unsigned(temp_4) | input_data);
    assign temp_6 = temp_1[1:0];
    assign temp_7 = (($unsigned(($unsigned(((input_data & temp_4) + temp_3)) * input_data)) * temp_6[2:2]) | temp_0);
    assign temp_8 = ($signed(((temp_1 ^ temp_3[19:16]) >> temp_7)) << input_data);
    assign temp_9 = temp_5;
    assign temp_10 = $unsigned(((($signed(($signed((temp_4 ^ temp_2)) & temp_8)) - (~temp_5)) | temp_2[10:5]) & temp_7));
    assign temp_11 = ($unsigned(input_data) * temp_7);
    assign temp_12 = $unsigned(temp_4);
    assign temp_13 = ($signed((($unsigned(temp_11) + temp_7) * temp_8)) & temp_10);
    assign temp_14 = $unsigned(((((temp_13 | temp_2) ^ temp_10) - temp_3) - temp_3));
    assign temp_15 = ($signed(temp_2) >> temp_14);
    assign temp_16 = (($unsigned((($unsigned(((temp_7 & temp_10) ^ temp_12)) ^ temp_2) & temp_5)) - temp_13[2:0]) * temp_4);
    assign temp_17 = $signed((temp_7 + temp_11));

    assign output_data = (($unsigned((($unsigned(temp_12[17:16]) & temp_10) & temp_12)) + temp_3) - temp_2);

endmodule