module top (
    input [2:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;

    assign temp_0 = ((((((input_data & input_data) & input_data) + input_data) + input_data) ^ input_data) + input_data);
    assign temp_1 = (((((((input_data | temp_0) - temp_0) ^ temp_0[24:11]) * temp_0) + temp_0[24:13]) & input_data) + temp_0[22:0]);
    assign temp_2 = ((temp_0 + temp_1) + 13'd2817);
    assign temp_3 = (((((((temp_0 - temp_2) * temp_0) ^ temp_0) ^ temp_2) & temp_2) * input_data) & input_data);
    assign temp_4 = (input_data - temp_3);
    assign temp_5 = ((((((temp_0 ^ temp_3) * temp_4) - input_data) | temp_1) ^ temp_4) | temp_2[8:0]);
    assign temp_6 = (((((temp_0 - temp_2) * temp_5) ^ temp_3[2:0]) ^ temp_0) - temp_0[24:0]);
    assign temp_7 = ($unsigned((((((($unsigned(temp_1) ^ temp_1[8:0]) >= temp_6) != temp_5) | temp_3) <= temp_4) > temp_0[24:12])) < temp_4);
    assign temp_8 = (input_data * temp_5);
    assign temp_9 = ((((((temp_2 ^ temp_0) - temp_4) * temp_4) & temp_7) | temp_5) - temp_8);
    assign temp_10 = ((($signed(temp_3[2:1]) + temp_9) - temp_0) << temp_6);

    assign output_data = ((((((temp_10[29:3] & temp_5) * temp_4) ^ temp_3) & temp_2) * temp_8) | temp_5);

endmodule