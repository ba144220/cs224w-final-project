module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;

    assign temp_0 = $signed(input_data);
    assign temp_1 = $unsigned((($unsigned(($signed((($signed(input_data) - 26'd40298301) * input_data)) & temp_0)) | (~input_data)) - input_data));
    assign temp_2 = $signed(input_data);
    assign temp_3 = (input_data * temp_0);
    assign temp_4 = (((((($signed((input_data * temp_1)) & input_data) | -6'd16) + temp_2) - temp_3) - temp_0) & -6'd30);
    assign temp_5 = $unsigned(temp_4);
    assign temp_6 = $unsigned(((($unsigned(((($unsigned(input_data[2:1]) & temp_2) * 2'd3) & temp_0[6:5])) & input_data[1:0]) | (~input_data[3:2])) ^ (~temp_3)));
    assign temp_7 = $signed(((((($unsigned(temp_3) & temp_3) * temp_3) - temp_6[1:1]) ^ (~temp_3)) - temp_2[30:26]));
    assign temp_8 = $unsigned((($unsigned(temp_5) | temp_7) ^ temp_6[1:1]));
    assign temp_9 = (temp_5 + temp_8);
    assign temp_10 = ($signed(((((((temp_1 ^ temp_4) & temp_4) & input_data) & temp_0) * temp_6[1:1]) ^ input_data)) & temp_7);
    assign temp_11 = (($unsigned(((temp_3 - temp_10) == temp_2)) != input_data) - temp_2);
    assign temp_12 = (((($unsigned(((temp_4[5:2] + temp_0) - temp_7)) & temp_2) * (~input_data)) ^ temp_9) ^ temp_1);
    assign temp_13 = $unsigned(((($signed(((temp_8 - temp_10) + temp_8[18:8])) + temp_0[6:0]) ^ temp_4) & input_data));
    assign temp_14 = (((($signed(((($signed(temp_12) & temp_9) ^ temp_2) | temp_3)) + temp_0) + temp_5) + temp_2) ^ temp_0);

    assign output_data = ($unsigned(((temp_2 + temp_10) - temp_13[11:8])) ^ temp_5);

endmodule