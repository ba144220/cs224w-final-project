module top (
    input [11:0] input_data,
    output [8:0] output_data
);

    logic [22:0] temp_0;
    logic [1:0] temp_1;
    logic [29:0] temp_2;
    logic [15:0] temp_3;
    logic [3:0] temp_4;
    logic [10:0] temp_5;
    logic [7:0] temp_6;
    logic [23:0] temp_7;
    logic [30:0] temp_8;
    logic [15:0] temp_9;
    logic [24:0] temp_10;
    logic [6:0] temp_11;
    logic [15:0] temp_12;
    logic [0:0] temp_13;
    logic [13:0] temp_14;
    logic [26:0] temp_15;
    logic [17:0] temp_16;

    assign temp_0 = (((input_data * input_data) * input_data) == input_data);
    assign temp_1 = $unsigned(($unsigned((temp_0 + temp_0)) - temp_0));
    assign temp_2 = temp_0;
    assign temp_3 = ($unsigned((((temp_1[1:1] - temp_2[29:9]) * temp_1[1:1]) & (~temp_0))) ^ (~temp_1));
    assign temp_4 = ($signed((((temp_0 + input_data[10:7]) - input_data[10:7]) * temp_3[15:14])) ^ input_data[5:2]);
    assign temp_5 = ((temp_2 & temp_2) & temp_2);
    assign temp_6 = $unsigned(((temp_1 * input_data[11:4]) * input_data[7:0]));
    assign temp_7 = $unsigned((((temp_2[29:6] | temp_5) & input_data) & (~temp_0)));
    assign temp_8 = $signed(((temp_5 * (~temp_5)) & temp_5));
    assign temp_9 = input_data;
    assign temp_10 = {12'b0, (((temp_6 - (~temp_4)) * temp_4[3:3]) * temp_2[29:18])};
    assign temp_11 = (temp_7 ^ temp_0);
    assign temp_12 = ((temp_0 + temp_8) ^ temp_10);
    assign temp_13 = $signed(($signed(((temp_11 >> temp_2) * (~temp_8[30:8]))) - temp_0));
    assign temp_14 = temp_7;
    assign temp_15 = temp_4;
    assign temp_16 = $signed((((temp_11 + temp_9) <= temp_7) <= (~temp_7)));

    assign output_data = temp_12;

endmodule