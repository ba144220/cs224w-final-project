module top (
    input [5:0] input_data,
    output [9:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;

    assign temp_0 = (($signed(input_data) - input_data) & input_data);
    assign temp_1 = ($signed(($signed(temp_0) | temp_0)) + input_data);
    assign temp_2 = ($signed((($unsigned(($signed(($unsigned(($unsigned((($unsigned(($unsigned(($unsigned(temp_0) & temp_0)) + temp_0)) - input_data) & temp_1[2:0])) * input_data)) | input_data)) * temp_1)) + temp_0[6:0]) ^ (~temp_1[2:0]))) * temp_1);
    assign temp_3 = $signed(($unsigned(temp_2[17:0]) & temp_1));
    assign temp_4 = ($unsigned(($unsigned(temp_3) + temp_1)) == temp_2);
    assign temp_5 = $signed(($unsigned(($signed(($signed(($unsigned((($signed(($signed((($signed(temp_0) | input_data) ^ temp_2)) * temp_1[23:0])) & (~temp_0)) | temp_4)) + temp_1[4:0])) - 31'd1719179043)) | temp_0)) + temp_3));
    assign temp_6 = ((($signed((($unsigned(temp_1) & temp_4) + temp_3[4:0])) ^ temp_0) & temp_0) * temp_5[27:0]);
    assign temp_7 = temp_4 ? temp_4 : temp_0;
    assign temp_8 = temp_3[1:0];
    assign temp_9 = $signed((($unsigned(($unsigned(($unsigned(($unsigned((($unsigned(((input_data >= temp_6) - temp_3)) != temp_8) > temp_8)) << temp_8)) != temp_4)) >= temp_5)) & temp_8[12:0]) + temp_3));
    assign temp_10 = ($signed((temp_4 * temp_1[9:0])) ^ temp_5[11:0]);
    assign temp_11 = ($signed(($unsigned(temp_10) | temp_5)) | temp_5);
    assign temp_12 = $unsigned((($unsigned(temp_5) + temp_8[6:0]) * temp_7));

    assign output_data = (temp_2[17:0] * temp_3);

endmodule