module top (
    input [4:0] input_data,
    output [9:0] output_data
);

    logic [25:0] temp_0;
    logic [3:0] temp_1;
    logic [4:0] temp_2;
    logic [6:0] temp_3;
    logic [23:0] temp_4;
    logic [3:0] temp_5;
    logic [13:0] temp_6;
    logic [2:0] temp_7;
    logic [5:0] temp_8;
    logic [27:0] temp_9;
    logic [26:0] temp_10;
    logic [4:0] temp_11;
    logic [15:0] temp_12;
    logic [5:0] temp_13;
    logic [27:0] temp_14;

    assign temp_0 = ((((input_data | (~input_data)) - input_data) | input_data) - input_data);
    assign temp_1 = $signed((((temp_0 | temp_0) + (~temp_0)) ^ temp_0));
    assign temp_2 = {1'b0, temp_1};
    assign temp_3 = $signed((temp_1[1:0] & temp_1[2:0]));
    assign temp_4 = {13'b0, ((temp_0[8:0] ^ (~temp_3)) | temp_2)};
    assign temp_5 = ((((((temp_3 ^ (~temp_1[1:0])) | temp_0) + input_data[3:0]) | temp_0[16:0]) & temp_1[2:0]) ^ temp_0);
    assign temp_6 = (((((temp_2 - temp_4) - temp_3) + input_data) * temp_5) - temp_2);
    assign temp_7 = $unsigned(temp_5);
    assign temp_8 = (((((input_data - temp_7) ^ input_data) ^ temp_2) * temp_3) + input_data);
    assign temp_9 = (temp_7 - temp_7);
    assign temp_10 = $signed(((((temp_1 - temp_9) <= temp_7) | (~input_data)) - temp_5[1:0]));
    assign temp_11 = (((((temp_7 & temp_2) | (~temp_6)) | temp_0) + input_data) - temp_2);
    assign temp_12 = $signed((((temp_11[1:0] * temp_10[9:0]) + temp_1) * temp_0));
    assign temp_13 = $unsigned(((((((temp_4[23:9] + temp_11) & temp_10) | temp_3) ^ temp_5) * temp_0[13:0]) * temp_11));
    assign temp_14 = (temp_2[4:0] - (~temp_8));

    assign output_data = (((temp_3[5:0] * temp_10) != temp_7[1:0]) <= temp_10);

endmodule