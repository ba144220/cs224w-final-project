module top (
    input [2:0] input_data,
    output [2:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;
    logic [17:0] temp_12;
    logic [2:0] temp_13;
    logic [1:0] temp_14;

    assign temp_0 = (((((input_data | input_data) - input_data) - input_data) * input_data) & input_data);
    assign temp_1 = $unsigned(((((((((input_data * input_data) * input_data) * input_data) | temp_0) ^ (~temp_0)) | temp_0) ^ (~24'd8371887)) + temp_0[5:2]));
    assign temp_2 = $signed(input_data);
    assign temp_3 = input_data;
    assign temp_4 = (input_data & temp_1);
    assign temp_5 = temp_3;
    assign temp_6 = (((temp_1 ^ temp_3) * temp_5[13:1]) & temp_5);
    assign temp_7 = ((((((temp_3 - temp_3) | (~temp_2)) & (~input_data)) >> temp_4[16:1]) - temp_3) ^ temp_0[5:5]);
    assign temp_8 = temp_0 ? (((((temp_7 ^ (~input_data)) | temp_6) | temp_5) + input_data) - temp_5) : $unsigned((temp_2 ^ temp_5));
    assign temp_9 = ((((((((temp_6 | temp_1) & input_data) & temp_1) - input_data) | temp_2) - temp_3) | input_data) & temp_8);
    assign temp_10 = ((((input_data & temp_7[10:5]) * temp_6) - temp_8) * (~temp_4));
    assign temp_11 = $unsigned(((temp_3 | temp_1) * temp_5[13:8]));
    assign temp_12 = $unsigned(((((temp_3 * temp_2) ^ temp_11) << temp_11) - temp_6));
    assign temp_13 = temp_11;
    assign temp_14 = $signed(((((((temp_5 + temp_12) * temp_11) | (~temp_2[10:8])) | temp_1) + temp_7) + temp_8));

    assign output_data = (((((((temp_14 * temp_1) ^ temp_3[19:3]) >> (~temp_0)) + temp_2) + temp_13) ^ temp_7) + temp_9);

endmodule