module top (
    input [5:0] input_data,
    output [2:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;

    assign temp_0 = (((((((((((input_data - input_data) + (~input_data)) * input_data) & input_data) * 9'd222) ^ input_data) * input_data) ^ input_data) ^ input_data) | input_data) * input_data);
    assign temp_1 = 1'd1 ? $signed((temp_0 | temp_0[8:1])) : (((((input_data | temp_0) ^ temp_0) & input_data) + temp_0) ^ temp_0[8:6]);
    assign temp_2 = $signed((((((temp_1[1:0] | temp_0) - temp_0[6:0]) - temp_0[4:0]) - temp_0) - input_data));
    logic [34:0] expr_957438;
    assign expr_957438 = (((((temp_0[8:1] & input_data[5:1]) ^ temp_2) | (~temp_0)) - temp_2) + (~temp_2));
    assign temp_3 = expr_957438[4:0];
    assign temp_4 = (((((temp_0 | temp_0) + temp_3[3:0]) | temp_3) + temp_0[8:2]) - temp_2);
    assign temp_5 = temp_3 ? $unsigned(temp_3[4:4]) : ($signed(((((temp_1 | temp_3[4:1]) | temp_2) | temp_0) + temp_1[23:3])) & temp_0);
    assign temp_6 = (temp_5 - (~temp_0));
    logic [36:0] expr_979135;
    assign expr_979135 = (((((((((((temp_3 + temp_1) ^ temp_4) - temp_3) ^ temp_1) - temp_4) | temp_2) - temp_2) ^ temp_4) + temp_5[13:0]) + (~temp_1)) - temp_1);
    assign temp_7 = expr_979135[14:0];

    assign output_data = temp_1[9:0];

endmodule