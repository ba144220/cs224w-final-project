module top (
    input [11:0] input_data,
    output [16:0] output_data
);

    logic [22:0] temp_0;
    logic [1:0] temp_1;
    logic [29:0] temp_2;
    logic [15:0] temp_3;
    logic [3:0] temp_4;
    logic [10:0] temp_5;
    logic [7:0] temp_6;
    logic [23:0] temp_7;
    logic [30:0] temp_8;
    logic [15:0] temp_9;
    logic [24:0] temp_10;
    logic [6:0] temp_11;
    logic [15:0] temp_12;

    assign temp_0 = input_data[4:4] ? ($unsigned(23'd2328130) | (~input_data)) : (input_data - input_data);
    assign temp_1 = (input_data[10:9] ^ temp_0);
    assign temp_2 = {28'b0, $signed(temp_1)};
    assign temp_3 = {15'b0, (input_data <= (~temp_1[1:0]))};
    assign temp_4 = $signed(((($unsigned((temp_0 - temp_1)) + input_data[9:6]) * temp_3[15:0]) * 4'd4));
    assign temp_5 = $signed(((temp_1 & temp_2) & temp_4));
    assign temp_6 = ((temp_4 ^ temp_5) | (~input_data[8:1]));
    assign temp_7 = (($signed((temp_2 ^ input_data)) * input_data) * temp_5);
    assign temp_8 = (($unsigned(((temp_0 | temp_3) - temp_2[6:0])) & temp_6) * temp_4);
    assign temp_9 = ($signed(($signed(temp_5) | temp_5)) - temp_5);
    assign temp_10 = ($signed(($signed(((temp_4 & input_data) * temp_5)) + temp_9)) & temp_4);
    assign temp_11 = ((($signed(temp_1[1:0]) * temp_5) | temp_0) | temp_6);
    assign temp_12 = ($signed(((temp_4 * temp_11) * temp_7)) & (~temp_0[8:0]));

    assign output_data = temp_0[4:0];

endmodule