module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;

    assign temp_0 = {1'b0, $signed(((input_data + input_data) & input_data))};
    assign temp_1 = ((input_data | temp_0) | temp_0);
    assign temp_2 = ((temp_0 - input_data) ^ input_data);
    assign temp_3 = temp_0[5:5];
    assign temp_4 = {16'b0, temp_1[23:23]};
    assign temp_5 = 14'd692;
    assign temp_6 = input_data[2:2] ? (($signed(temp_1[23:12]) >= temp_5) != temp_2) : ($unsigned(temp_1) >> temp_1);
    assign temp_7 = ($unsigned(temp_5) != temp_1);
    assign temp_8 = ($signed(temp_6) ^ temp_1);
    assign temp_9 = temp_6[2:1];

    assign output_data = temp_0;

endmodule