module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;

    assign temp_0 = $signed(input_data);
    assign temp_1 = $signed((input_data - temp_0));
    assign temp_2 = ($signed(($signed(temp_1) + temp_1)) ^ temp_1);
    assign temp_3 = ($unsigned(temp_2) ^ input_data);
    logic [9:0] expr_647736;
    assign expr_647736 = temp_3;
    assign temp_4 = expr_647736[5:0];
    assign temp_5 = $signed(($signed(temp_1[25:2]) & temp_2));
    assign temp_6 = temp_2;
    assign temp_7 = temp_0;
    assign temp_8 = $signed(temp_3);
    assign temp_9 = input_data[5:2];
    assign temp_10 = temp_2;
    assign temp_11 = $unsigned(($signed(($unsigned(temp_5) + (~temp_4))) * temp_0));
    logic [21:0] expr_83560;
    assign expr_83560 = ($unsigned((temp_6 - temp_9)) | temp_1[20:0]);
    assign temp_12 = expr_83560[17:0];
    assign temp_13 = ((temp_1 & temp_4) + temp_9);
    assign temp_14 = temp_1;
    assign temp_15 = $signed(($unsigned(17'd81740) + temp_7));
    assign temp_16 = temp_14;

    assign output_data = ((temp_11 & temp_2) * (~temp_6));

endmodule