module top (
    input [2:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;

    assign temp_0 = {19'b0, ($unsigned(($unsigned(($unsigned(input_data) ^ input_data)) ^ input_data)) + input_data)};
    assign temp_1 = input_data[0:0] ? ($signed(($unsigned(input_data) | temp_0)) ^ input_data) : ($signed(($unsigned(($unsigned(temp_0) & temp_0)) - input_data)) - input_data);
    assign temp_2 = temp_0 ? ($unsigned(($signed(input_data) - temp_0)) * temp_1) : $signed(($unsigned(($signed(temp_0) & input_data)) & input_data));
    assign temp_3 = temp_1;
    assign temp_4 = $signed(($unsigned((($signed(temp_1[5:0]) + input_data) ^ temp_2)) * input_data));
    assign temp_5 = ((($signed((($unsigned(temp_3) | input_data) + temp_2)) ^ temp_2) | temp_1) ^ temp_4);
    assign temp_6 = temp_5 ? $signed((16'd11004 - temp_2[12:4])) : ($unsigned(($signed(($signed(($unsigned(($unsigned(input_data) - temp_3)) - temp_1[1:0])) - temp_2)) + input_data)) - 16'd37662);
    assign temp_7 = $unsigned(($unsigned(($signed(($unsigned(($signed(($signed(($signed(($unsigned(input_data) ^ input_data)) | temp_1)) * (~temp_0))) - 14'd14710)) & temp_4[5:5])) * temp_2)) * (~input_data)));
    assign temp_8 = temp_7;
    assign temp_9 = $unsigned(((($unsigned(($unsigned(input_data[2:1]) & temp_1)) * temp_7) - temp_0[22:0]) ^ temp_3[2:2]));
    assign temp_10 = {15'b0, $signed(($unsigned(($unsigned(($unsigned(($unsigned(temp_5[8:4]) + input_data)) << input_data)) ^ input_data)) + temp_7))};
    assign temp_11 = ($signed(((temp_7 - temp_1) & temp_9)) - temp_5);
    assign temp_12 = ($unsigned(($signed((($unsigned(temp_10) + temp_6) & temp_0)) - temp_0)) | temp_2[8:0]);
    assign temp_13 = ($unsigned(($unsigned(($signed((($signed((temp_7 + temp_7)) ^ temp_12) - temp_9)) ^ temp_8)) * temp_0)) ^ temp_7);

    assign output_data = ($signed(temp_11) ^ temp_3);

endmodule