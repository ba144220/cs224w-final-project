module top (
    input [2:0] input_data,
    output [4:0] output_data
);

    logic [23:0] temp_0;
    logic [30:0] temp_1;
    logic [4:0] temp_2;
    logic [0:0] temp_3;
    logic [30:0] temp_4;
    logic [16:0] temp_5;
    logic [14:0] temp_6;

    assign temp_0 = (($signed(($signed(((($signed((input_data - input_data)) + input_data) & input_data) & input_data)) * input_data)) ^ input_data) | input_data);
    assign temp_1 = ($unsigned(($signed(($signed(($unsigned(($unsigned((($unsigned((((temp_0 | temp_0[21:0]) + temp_0[14:0]) + input_data)) * temp_0[23:20]) * input_data)) * input_data)) | input_data)) * temp_0)) + temp_0[21:0])) | (~input_data));
    assign temp_2 = ($unsigned(($unsigned(($unsigned(($signed(($signed(($unsigned(($unsigned(($unsigned(($unsigned(temp_1) & temp_0)) * temp_0)) ^ input_data)) | temp_0[23:7])) * temp_0)) * temp_1)) & input_data)) + input_data)) | input_data);
    assign temp_3 = (($signed((($signed(($signed(($unsigned((($unsigned(($signed(temp_2) <= temp_0)) > input_data[0:0]) * (~temp_1))) == temp_1[9:0])) + temp_0)) + input_data[2:2]) < temp_2)) * temp_2) == input_data[0:0]);
    assign temp_4 = (($unsigned(($unsigned((($signed(temp_1) | temp_3) | temp_2)) | (~temp_0))) - temp_3) + temp_0[4:0]);
    assign temp_5 = $unsigned(temp_1[24:0]);
    assign temp_6 = $signed(($unsigned(($signed(temp_1) & temp_4)) & temp_1));

    assign output_data = $signed(((($unsigned(($unsigned(($signed((($signed(temp_4) - temp_1) ^ temp_4)) | temp_4)) - temp_1)) ^ temp_3) + temp_3) + temp_3));

endmodule