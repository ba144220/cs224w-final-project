module top (
    input [3:0] input_data,
    output [4:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;
    logic [16:0] temp_6;
    logic [14:0] temp_7;
    logic [12:0] temp_8;
    logic [30:0] temp_9;
    logic [30:0] temp_10;
    logic [25:0] temp_11;
    logic [9:0] temp_12;
    logic [14:0] temp_13;

    assign temp_0 = ((((input_data + input_data) << input_data) >> (~input_data)) * input_data);
    assign temp_1 = {12'b0, $unsigned((((temp_0 + input_data) | input_data) * temp_0))};
    assign temp_2 = (((31'd1421437244 | temp_0[8:1]) | input_data) ^ input_data);
    assign temp_3 = temp_1;
    assign temp_4 = ((temp_2[20:0] * temp_2) >> temp_0[8:6]);
    assign temp_5 = ((temp_3 | input_data) * temp_3[4:3]);
    assign temp_6 = {13'b0, input_data};
    assign temp_7 = ((temp_2 + input_data) * temp_5);
    assign temp_8 = ((((input_data + temp_4) * temp_3[2:0]) | temp_7) | temp_0);
    assign temp_9 = ((input_data * input_data) & (~temp_4));
    assign temp_10 = (temp_0[8:8] ^ temp_1);
    assign temp_11 = ((((temp_9 >= temp_8) ^ temp_5) <= temp_9[14:0]) + input_data);
    assign temp_12 = ((((temp_9 ^ temp_2) ^ (~temp_2)) + (~temp_11)) | temp_11);
    assign temp_13 = temp_9;

    assign output_data = ((((temp_8 ^ temp_2) ^ temp_7) & temp_11) - temp_2);

endmodule