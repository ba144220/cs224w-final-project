module top (
    input [2:0] input_data,
    output [31:0] output_data
);

    logic [16:0] temp_0;
    logic [2:0] temp_1;
    logic [0:0] temp_2;
    logic [9:0] temp_3;
    logic [30:0] temp_4;
    logic [23:0] temp_5;
    logic [20:0] temp_6;

    assign temp_0 = ((((input_data - input_data) + input_data) & input_data) ^ input_data);
    assign temp_1 = (((((((temp_0 & temp_0[7:0]) * input_data) ^ temp_0) | temp_0) + temp_0[15:0]) | temp_0) & temp_0);
    assign temp_2 = temp_1 ? ((((temp_1 & temp_1) ^ input_data[2:2]) | temp_1) * temp_1) : $signed((((((((temp_1 >> temp_0) ^ temp_0) - temp_0) | input_data[1:1]) * input_data[1:1]) | temp_0) + temp_1));
    assign temp_3 = $unsigned(((((((((temp_0[7:0] ^ temp_0) ^ temp_0) ^ temp_1) - temp_2) - temp_0) & temp_0) ^ temp_2) - temp_0));
    assign temp_4 = {30'b0, temp_2};
    assign temp_5 = (((((((input_data == input_data) == temp_1) != temp_2) ^ temp_1) < temp_0) > temp_0) <= temp_3);
    assign temp_6 = $signed(temp_4);

    assign output_data = $unsigned((((((((temp_5 - temp_6) + temp_2) ^ temp_2) | temp_6) - temp_4) * temp_2) + temp_2));

endmodule