module top (
    input [5:0] input_data,
    output [9:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;

    logic [11:0] expr_319932;
    assign expr_319932 = (((($unsigned(($signed(7'd6) ^ input_data)) ^ input_data) | (~input_data)) | input_data) * input_data);
    assign temp_0 = expr_319932[6:0];
    assign temp_1 = input_data;
    assign temp_2 = ($signed(temp_1) | temp_0);
    assign temp_3 = $unsigned(((temp_0 ^ temp_1) - temp_0));
    assign temp_4 = (((((temp_0 - (~temp_0)) + temp_1[25:17]) ^ input_data) - (~temp_1)) + temp_1);
    assign temp_5 = (input_data[4:0] & temp_3);
    assign temp_6 = (($unsigned((((((((($unsigned(temp_5) & (~2'd1)) * temp_0) & (~input_data[1:0])) | 2'd3) - temp_4) | temp_0) | (~temp_0)) * temp_0)) & temp_3) * temp_3);
    assign temp_7 = $unsigned(($signed((((((($signed(temp_6) * temp_2) + temp_3) & (~temp_2)) + temp_2) | temp_4) ^ (~temp_3))) * temp_6));
    logic [25:0] expr_612545;
    assign expr_612545 = temp_1;
    assign temp_8 = expr_612545[18:0];
    assign temp_9 = ((($signed((((((((temp_1 ^ temp_4) & temp_4) & temp_6) | temp_2) & temp_0) * temp_4) & temp_1)) - temp_8) - temp_5) | temp_2);
    logic [31:0] expr_338007;
    assign expr_338007 = $unsigned(((((((((temp_4 - temp_4) - temp_6) - temp_1) & temp_8) ^ (~temp_6)) & temp_5) + temp_3) & temp_5));
    assign temp_10 = expr_338007[14:0];

    assign output_data = $signed((($signed((((temp_0 | temp_3) - temp_4) + (~temp_1))) ^ temp_0[6:0]) ^ temp_5));

endmodule