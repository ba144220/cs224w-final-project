module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;

    assign temp_0 = input_data;
    assign temp_1 = ($signed(temp_0) - input_data);
    assign temp_2 = {4'b0, (temp_1 + (~temp_1))};
    assign temp_3 = (($unsigned(temp_2) - -10'd118) + temp_0[6:3]);
    assign temp_4 = temp_3;
    assign temp_5 = (temp_1[25:2] & temp_2);
    assign temp_6 = temp_4[5:1] ? ($signed((2'd3 ^ input_data[2:1])) - (~temp_1)) : temp_2;
    assign temp_7 = ((temp_1 - temp_5) - temp_5);
    assign temp_8 = temp_4[5:2];
    assign temp_9 = (temp_2[29:0] * temp_6);
    assign temp_10 = $unsigned((temp_9 * temp_2[3:0]));
    assign temp_11 = temp_6 ? ($unsigned(24'd12276977) | input_data) : ($signed(temp_2[30:16]) ^ temp_0[6:3]);
    assign temp_12 = (temp_10[1:0] | temp_8);
    assign temp_13 = (temp_10 | temp_12);
    assign temp_14 = temp_10[14:1];
    assign temp_15 = temp_2;
    assign temp_16 = temp_3 ? ((temp_12 & temp_9) & temp_12) : $unsigned(((temp_12 - temp_14) * temp_8));

    assign output_data = temp_1 ? $unsigned(($signed(($signed(temp_8[8:0]) - temp_3)) ^ temp_9)) : ($unsigned(temp_4[5:3]) & temp_16[3:0]);

endmodule