module top (
    input [2:0] input_data,
    output [11:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;

    assign temp_0 = (($unsigned(((($unsigned(((input_data + input_data) & input_data)) + input_data) + input_data) - input_data)) + input_data) | input_data);
    assign temp_1 = $unsigned(($signed(($signed(($unsigned(($signed((input_data * temp_0[24:17])) * temp_0)) ^ input_data)) + temp_0[24:13])) - temp_0[24:3]));
    assign temp_2 = ($unsigned(((($signed(($unsigned((($unsigned(temp_0) ^ temp_1) | temp_0)) | temp_1)) ^ temp_0) - temp_0) + input_data)) | temp_0);
    assign temp_3 = (((((temp_1 ^ temp_2) * temp_0) * temp_1) ^ temp_2) | temp_0[24:24]);
    assign temp_4 = ($unsigned(($signed((($unsigned(temp_3) - input_data) - temp_0)) & input_data)) + temp_2[12:10]);
    assign temp_5 = $signed(($signed(($unsigned(input_data) | temp_1)) ^ temp_3));
    assign temp_6 = (($signed((temp_5 ^ temp_1)) * input_data) >> temp_3);
    assign temp_7 = $unsigned((($signed(($unsigned((($signed(($signed((temp_1 & temp_6)) | temp_1)) * temp_0) - temp_0)) & temp_4[5:5])) * temp_2) * temp_6));
    assign temp_8 = temp_7;

    assign output_data = ($signed((($unsigned(($unsigned(temp_4) & temp_1)) * temp_7) - temp_8[25:22])) ^ temp_6);

endmodule