module top (
    input [5:0] input_data,
    output [37:0] output_data
);

    logic [8:0] temp_0;
    logic [23:0] temp_1;
    logic [30:0] temp_2;
    logic [4:0] temp_3;
    logic [0:0] temp_4;
    logic [30:0] temp_5;

    assign temp_0 = (($unsigned(($signed(input_data) & input_data)) & (~input_data)) + input_data);
    assign temp_1 = $unsigned(((((((temp_0 - temp_0) | input_data) ^ 24'd5472715) | input_data) * temp_0) + temp_0[7:0]));
    assign temp_2 = $unsigned((($signed(((($signed(temp_0) + temp_0) * temp_0) ^ input_data)) | temp_0) & input_data));
    assign temp_3 = (($signed(($signed((($unsigned(temp_2[22:0]) + input_data[5:1]) - (~temp_1))) + input_data[4:0])) - temp_2) - temp_0[4:0]);
    assign temp_4 = (($signed((temp_2 + temp_2)) & temp_3) & input_data[4:4]);
    assign temp_5 = ($signed((((temp_4 - temp_4) + temp_0) & temp_4)) + temp_1);

    assign output_data = $signed(((($signed(($signed(($signed((($unsigned(temp_0) | temp_4) - temp_0)) + temp_4)) | temp_2)) ^ temp_5) | (~temp_3)) ^ temp_3));

endmodule