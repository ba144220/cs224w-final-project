module top (
    input [2:0] input_data,
    output [23:0] output_data
);

    logic [24:0] temp_0;
    logic [8:0] temp_1;
    logic [12:0] temp_2;
    logic [2:0] temp_3;
    logic [5:0] temp_4;
    logic [8:0] temp_5;
    logic [15:0] temp_6;
    logic [13:0] temp_7;
    logic [25:0] temp_8;
    logic [1:0] temp_9;
    logic [29:0] temp_10;
    logic [31:0] temp_11;
    logic [29:0] temp_12;
    logic [24:0] temp_13;
    logic [31:0] temp_14;

    assign temp_0 = (((25'd27357858 > input_data) - input_data) - (~input_data));
    assign temp_1 = (temp_0 & input_data);
    assign temp_2 = ((input_data * temp_1[8:4]) * temp_1[5:0]);
    logic [12:0] expr_73374;
    assign expr_73374 = (temp_0[24:13] * input_data);
    assign temp_3 = expr_73374[2:0];
    assign temp_4 = input_data;
    assign temp_5 = temp_4;
    logic [27:0] expr_221475;
    assign expr_221475 = $signed((((temp_4 & temp_0) & temp_4) + input_data));
    assign temp_6 = expr_221475[15:0];
    assign temp_7 = temp_5;
    assign temp_8 = (((temp_4 & temp_4[4:0]) ^ input_data) + temp_5);
    assign temp_9 = ((temp_6 | input_data[1:0]) & input_data[2:1]);
    assign temp_10 = (((temp_8 | temp_3) ^ temp_9) | temp_4[4:0]);
    assign temp_11 = ((temp_0[24:5] ^ temp_1) * temp_5[2:0]);
    assign temp_12 = (temp_3[1:0] * temp_1[8:3]);
    assign temp_13 = (((temp_2[12:6] & temp_2) == temp_6) ^ temp_11);
    assign temp_14 = (temp_8 * temp_9);

    logic [32:0] expr_243915;
    assign expr_243915 = (temp_14 * temp_11[31:5]);
    assign output_data = temp_5 ? (((temp_2[12:3] & temp_9) | temp_14) ^ temp_5) : expr_243915[23:0];

endmodule