module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;

    assign temp_0 = $signed(input_data);
    assign temp_1 = ($signed(($signed(temp_0) - input_data)) | input_data);
    assign temp_2 = temp_1;
    assign temp_3 = ($signed(($signed(($signed(($signed((temp_2 - input_data)) | temp_0)) + input_data)) ^ temp_2[30:20])) & temp_0[6:1]);
    assign temp_4 = ($unsigned(temp_0) - temp_3);
    assign temp_5 = ($signed(temp_3) & temp_3[9:5]);
    assign temp_6 = input_data[4:4] ? ($unsigned(((input_data[1:0] & temp_3) * temp_3)) ^ temp_2) : (($unsigned((input_data[1:0] - temp_3)) + temp_1[9:0]) - temp_1);
    assign temp_7 = $signed(temp_6);
    assign temp_8 = ($unsigned(($unsigned(temp_7) * temp_7)) * temp_6);
    assign temp_9 = temp_2;
    assign temp_10 = temp_8;
    assign temp_11 = (($unsigned((temp_10[1:0] | temp_8)) | temp_9) * temp_1);
    assign temp_12 = (((($unsigned((temp_2 * (~temp_0))) ^ temp_1) - temp_7) | temp_11) | temp_11);
    logic [20:0] expr_968884;
    assign expr_968884 = ($unsigned(($unsigned(temp_8) * temp_6)) * temp_4);
    assign temp_13 = expr_968884[11:0];
    assign temp_14 = ((temp_9 | (~temp_3[9:1])) | temp_10);

    assign output_data = (($unsigned(($unsigned((($signed(temp_0) <= temp_6) | temp_8)) < temp_0[6:6])) * temp_1) != temp_8);

endmodule