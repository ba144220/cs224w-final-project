module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;
    logic [13:0] temp_16;
    logic [1:0] temp_17;

    assign temp_0 = ($unsigned((input_data + input_data)) - input_data);
    assign temp_1 = ((temp_0 * temp_0[4:0]) | input_data);
    assign temp_2 = ((input_data * temp_0) + temp_0[6:3]);
    assign temp_3 = temp_2;
    logic [31:0] expr_65231;
    assign expr_65231 = (temp_1[25:2] & temp_2);
    assign temp_4 = expr_65231[5:0];
    assign temp_5 = temp_1 ? (input_data ^ input_data) : (((input_data + temp_1) * temp_2) ^ input_data);
    assign temp_6 = (input_data[2:1] | temp_5);
    assign temp_7 = (temp_2[30:6] != temp_4);
    assign temp_8 = ((input_data & temp_5) > temp_0);
    assign temp_9 = input_data[2:2] ? (($unsigned(temp_6) & temp_7) * temp_6) : (((temp_2 & (~input_data)) * temp_1) - temp_4);
    assign temp_10 = (($unsigned((input_data | temp_6)) - temp_9) | temp_9);
    assign temp_11 = temp_1;
    assign temp_12 = (((temp_1 ^ temp_10) & temp_4) & input_data);
    assign temp_13 = (((temp_6 + temp_10) * temp_10) - temp_2);
    assign temp_14 = (temp_5[3:0] + temp_10);
    assign temp_15 = temp_8;
    assign temp_16 = (($unsigned(($unsigned(temp_12) & temp_12[1:0])) - temp_3) ^ temp_14);
    assign temp_17 = (temp_9 < temp_1);

    assign output_data = ((temp_7 ^ temp_1) + temp_5);

endmodule