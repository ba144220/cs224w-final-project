module top (
    input [2:0] input_data,
    output [5:0] output_data
);

    logic [5:0] temp_0;
    logic [23:0] temp_1;
    logic [10:0] temp_2;
    logic [19:0] temp_3;
    logic [16:0] temp_4;
    logic [13:0] temp_5;
    logic [2:0] temp_6;
    logic [10:0] temp_7;
    logic [27:0] temp_8;
    logic [25:0] temp_9;
    logic [23:0] temp_10;
    logic [28:0] temp_11;
    logic [17:0] temp_12;
    logic [2:0] temp_13;
    logic [1:0] temp_14;
    logic [23:0] temp_15;
    logic [29:0] temp_16;
    logic [20:0] temp_17;
    logic [24:0] temp_18;

    assign temp_0 = $unsigned((6'd17 | input_data));
    assign temp_1 = ($unsigned(($signed(temp_0) | temp_0)) & temp_0);
    assign temp_2 = {6'b0, ((input_data * input_data) + input_data)};
    assign temp_3 = ($signed(($signed(input_data) * temp_0[5:1])) + temp_0[1:0]);
    assign temp_4 = temp_1[23:12] ? temp_0 : ($signed(($signed(($signed(temp_0[2:0]) | temp_3)) & temp_1)) - temp_0);
    assign temp_5 = ($unsigned(($signed(temp_1[14:0]) - (~temp_0[5:2]))) ^ temp_2);
    assign temp_6 = temp_3 ? temp_0 : $signed(temp_1);
    logic [20:0] expr_84421;
    assign expr_84421 = $signed(($signed(temp_0) + temp_3));
    assign temp_7 = expr_84421[10:0];
    assign temp_8 = $signed(($signed(($signed(temp_0) + temp_7)) & temp_6));
    assign temp_9 = temp_6;
    assign temp_10 = $unsigned(temp_5);
    assign temp_11 = temp_2;
    assign temp_12 = (temp_6 | temp_4);
    logic [30:0] expr_855240;
    assign expr_855240 = ($unsigned(($signed(temp_11) & temp_6)) & temp_1[7:0]);
    assign temp_13 = expr_855240[2:0];
    assign temp_14 = $unsigned(($unsigned(temp_7[10:10]) ^ temp_4));
    assign temp_15 = temp_5;
    assign temp_16 = ($signed(($signed(temp_12) ^ temp_5)) & input_data);
    assign temp_17 = ($signed(($unsigned(temp_9) + temp_6)) * temp_14);
    assign temp_18 = $unsigned(($signed(($signed(temp_14) - temp_14)) & temp_11));

    assign output_data = $signed((($unsigned(temp_9) + temp_11) + temp_5));

endmodule