module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [23:0] temp_0;
    logic [17:0] temp_1;
    logic [8:0] temp_2;
    logic [11:0] temp_3;
    logic [0:0] temp_4;
    logic [21:0] temp_5;
    logic [29:0] temp_6;

    assign temp_0 = {17'b0, (input_data - input_data)};
    assign temp_1 = (($unsigned((($unsigned((((((input_data & temp_0) ^ (~input_data)) < input_data) - 18'd103636) + input_data)) <= input_data) * temp_0)) | input_data) & temp_0);
    assign temp_2 = ((($signed((($signed(((((temp_0 + temp_0) * temp_0) ^ input_data) & temp_1)) + (~temp_0)) & temp_1[17:12])) * temp_0) | input_data) | input_data);
    logic [25:0] expr_674035;
    assign expr_674035 = ((temp_0 | (~temp_0)) ^ temp_2);
    assign temp_3 = expr_674035[11:0];
    assign temp_4 = (($signed(($signed((temp_0 > input_data[5:5])) > temp_3[11:10])) >= temp_1) <= (~temp_0[23:3]));
    assign temp_5 = ((((((temp_2 - temp_1[17:3]) * temp_0) - temp_4) + temp_3) - temp_2[8:3]) & temp_2[8:6]);
    assign temp_6 = (((($unsigned((($unsigned(temp_3) & temp_2) ^ temp_1[17:15])) ^ temp_1) - temp_2) + temp_4) + temp_1);

    assign output_data = (($signed(temp_2) | temp_1) + temp_2);

endmodule