module top (
    input [5:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;

    assign temp_0 = input_data;
    assign temp_1 = input_data;
    assign temp_2 = (((((input_data - temp_0) + input_data) & temp_1) + temp_1) * temp_0);
    assign temp_3 = ($signed(((temp_0 & (~temp_0)) | input_data)) * input_data);
    assign temp_4 = $unsigned((($signed(temp_1) | (~temp_3)) * temp_1));
    assign temp_5 = ((($signed(temp_0) ^ input_data[5:1]) | temp_1) * temp_4);
    assign temp_6 = ((($unsigned(input_data[3:2]) ^ temp_5) * input_data[1:0]) ^ temp_0);
    assign temp_7 = (($signed((((((temp_1 - temp_2) | temp_1) & temp_3) * temp_1) * temp_6)) * temp_6) * temp_3);
    assign temp_8 = ($unsigned(((((((temp_2 & (~temp_4)) * (~temp_1)) - temp_4) ^ temp_5) | temp_7) * temp_1)) * temp_5);

    assign output_data = temp_1;

endmodule