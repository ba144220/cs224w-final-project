module top (
    input [4:0] input_data,
    output [16:0] output_data
);

    logic [22:0] temp_0;
    logic [1:0] temp_1;
    logic [29:0] temp_2;
    logic [15:0] temp_3;
    logic [3:0] temp_4;
    logic [10:0] temp_5;
    logic [7:0] temp_6;
    logic [23:0] temp_7;
    logic [30:0] temp_8;
    logic [15:0] temp_9;
    logic [24:0] temp_10;
    logic [6:0] temp_11;
    logic [15:0] temp_12;
    logic [0:0] temp_13;
    logic [13:0] temp_14;

    assign temp_0 = ($unsigned(23'd2328130) | (~input_data));
    assign temp_1 = ($signed(input_data[2:1]) - input_data[4:3]);
    assign temp_2 = ($unsigned(($unsigned(($unsigned((30'd657267987 & input_data)) + input_data)) | input_data)) - input_data);
    assign temp_3 = ($signed(($signed(16'd47530) * temp_2)) * input_data);
    assign temp_4 = ($signed(($signed(($unsigned(($unsigned(4'd1) & temp_1[1:0])) & temp_0)) | temp_3)) + temp_1);
    assign temp_5 = ($unsigned(($unsigned(input_data) & temp_2)) * temp_2);
    assign temp_6 = ($unsigned(($unsigned(input_data) ^ temp_4)) - input_data);
    assign temp_7 = ($unsigned(($unsigned(temp_3) * temp_0)) * temp_4[2:0]);
    assign temp_8 = ($signed(($unsigned(temp_1) + temp_4[3:0])) * input_data);
    assign temp_9 = temp_1;
    assign temp_10 = ($signed(($signed(((temp_4 & input_data) * temp_5)) + temp_9)) & temp_4);
    assign temp_11 = ($unsigned(($signed((input_data - (~temp_8))) * temp_9[1:0])) ^ temp_0);
    assign temp_12 = ($signed(($signed(($signed(temp_4) * temp_11)) - temp_8)) + temp_3[15:2]);
    assign temp_13 = temp_1[1:1];
    assign temp_14 = $signed(($signed(temp_9) ^ temp_1));

    assign output_data = ($unsigned((temp_0[10:0] - temp_9)) | temp_3);

endmodule