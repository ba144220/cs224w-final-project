module top (
    input [3:0] input_data,
    output [19:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;
    logic [16:0] temp_15;

    assign temp_0 = $signed(input_data);
    assign temp_1 = $signed((((((input_data & temp_0) + input_data) < temp_0) + temp_0) ^ temp_0[2:0]));
    assign temp_2 = (((temp_0 - temp_0[6:3]) * input_data) - input_data);
    assign temp_3 = ((temp_0 | temp_1) + input_data);
    assign temp_4 = input_data[3:3] ? (((($unsigned((((((($signed(temp_3) & temp_3) - input_data) * temp_3) + temp_0) - temp_3) ^ input_data)) + input_data) * 6'd59) & temp_0) & input_data) : (((($unsigned((input_data + temp_0)) * temp_0) - input_data) & temp_0) & input_data);
    assign temp_5 = $signed(($signed(input_data) * temp_2));
    assign temp_6 = ((((((((input_data[1:0] == temp_0) >= temp_4) >= temp_5) >= temp_2) - temp_1) >= temp_0) >= input_data[1:0]) - temp_3);
    assign temp_7 = ((((((($unsigned(((temp_2 ^ temp_3) * temp_4[2:0])) | temp_2) ^ input_data) & temp_3) * temp_0[5:0]) | temp_4) + temp_0) - input_data);
    assign temp_8 = ((((((((temp_4[5:2] - input_data) & temp_6[1:0]) * 19'd16123) & input_data) ^ input_data) + temp_5) + input_data) * 19'd331387);
    assign temp_9 = (((($signed((temp_8 - temp_1)) | input_data) + input_data) * temp_5) + temp_7);
    assign temp_10 = ((($unsigned((((temp_6 & input_data) * temp_1[9:0]) ^ temp_5[2:0])) * temp_7) + temp_1[11:0]) ^ temp_1);
    assign temp_11 = ((((temp_9 * temp_3[1:0]) + temp_4) & temp_6) != temp_0[6:2]);
    assign temp_12 = $unsigned(((((((((((temp_3 | temp_0[3:0]) | temp_0) & (~temp_5)) ^ temp_3[5:0]) + temp_10) | temp_10[7:0]) | temp_2) * temp_5) * temp_5[4:2]) - temp_1[21:0]));
    assign temp_13 = temp_1[25:20] ? (($signed(temp_7) ^ temp_4) + temp_8) : input_data;
    assign temp_14 = temp_0 ? ($signed(((($unsigned(((((temp_10[4:0] | temp_0[6:4]) | temp_5) | temp_0[3:0]) * temp_12[12:0])) | temp_7) * temp_10) - temp_5)) | temp_5) : (((((((temp_0[1:0] ^ temp_2) - (~temp_11)) - (~temp_0)) - input_data) * temp_12) | temp_6[1:0]) + temp_1[15:0]);
    assign temp_15 = $unsigned(((((temp_1 & temp_13[8:0]) - temp_9[2:0]) + temp_12) & temp_8));

    assign output_data = (((((temp_8 - temp_8) & temp_4) | temp_1) - temp_5) - temp_1[8:0]);

endmodule