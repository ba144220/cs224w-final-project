module top (
    input [3:0] input_data,
    output [9:0] output_data
);

    logic [6:0] temp_0;
    logic [25:0] temp_1;
    logic [30:0] temp_2;
    logic [9:0] temp_3;
    logic [5:0] temp_4;
    logic [4:0] temp_5;
    logic [1:0] temp_6;
    logic [25:0] temp_7;
    logic [18:0] temp_8;
    logic [3:0] temp_9;
    logic [14:0] temp_10;
    logic [23:0] temp_11;
    logic [17:0] temp_12;
    logic [11:0] temp_13;
    logic [6:0] temp_14;

    assign temp_0 = $signed(input_data);
    assign temp_1 = ($signed(($signed(temp_0) - input_data)) | input_data);
    assign temp_2 = {5'b0, temp_1};
    assign temp_3 = ($signed((($signed(($signed((temp_2 - input_data)) | temp_0[2:0])) + input_data) ^ temp_2)) * temp_1);
    assign temp_4 = ($signed(($signed(($signed(($signed(temp_1[2:0]) + temp_1)) <= temp_3)) & temp_1)) | temp_1);
    assign temp_5 = (($signed(($unsigned(($signed(($signed(temp_3) | input_data)) * input_data)) * input_data)) * temp_0) & temp_0);
    assign temp_6 = ($unsigned(temp_5) | temp_3);
    assign temp_7 = $unsigned(temp_0);
    assign temp_8 = ($signed((temp_6[1:0] | temp_5)) + temp_3);
    assign temp_9 = (($unsigned(temp_0[6:3]) + temp_7) * temp_2);
    assign temp_10 = $unsigned((($unsigned((($unsigned(temp_9) * temp_5) | temp_5)) + temp_2) | input_data));
    assign temp_11 = temp_10;
    assign temp_12 = $unsigned(($signed((($unsigned(((temp_11 ^ temp_10) * temp_6)) | temp_5) ^ temp_9)) ^ temp_9));
    assign temp_13 = ($unsigned(($signed(((temp_1 + temp_0) - temp_10)) * temp_11)) | temp_2);
    assign temp_14 = temp_4 ? (temp_0 > temp_8) : ($signed(($unsigned(($unsigned(temp_3[6:0]) * temp_13)) ^ temp_12)) * temp_10);

    assign output_data = temp_8 ? (temp_5 != temp_4[5:0]) : temp_0;

endmodule